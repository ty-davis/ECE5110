magic
tech sky130A
timestamp 1739990900
<< nwell >>
rect -2 197 215 488
<< nmos >>
rect 72 65 87 115
rect 108 65 123 115
<< pmos >>
rect 72 315 87 415
rect 126 315 141 415
<< ndiff >>
rect 36 107 72 115
rect 36 73 44 107
rect 61 73 72 107
rect 36 65 72 73
rect 87 65 108 115
rect 123 107 159 115
rect 123 73 134 107
rect 151 73 159 107
rect 123 65 159 73
<< pdiff >>
rect 36 407 72 415
rect 36 323 44 407
rect 61 323 72 407
rect 36 315 72 323
rect 87 315 126 415
rect 141 407 177 415
rect 141 323 152 407
rect 169 323 177 407
rect 141 315 177 323
<< ndiffc >>
rect 44 73 61 107
rect 134 73 151 107
<< pdiffc >>
rect 44 323 61 407
rect 152 323 169 407
<< psubdiff >>
rect 0 10 12 38
rect 201 10 213 38
<< nsubdiff >>
rect 16 442 28 470
rect 185 442 197 470
<< psubdiffcont >>
rect 12 10 201 38
<< nsubdiffcont >>
rect 28 442 185 470
<< poly >>
rect 72 415 87 428
rect 126 415 141 428
rect 72 301 87 315
rect 36 286 87 301
rect 36 252 52 286
rect 126 262 141 315
rect 19 244 52 252
rect 19 227 27 244
rect 44 227 52 244
rect 90 254 141 262
rect 90 237 98 254
rect 115 245 141 254
rect 115 237 123 245
rect 90 229 123 237
rect 19 219 52 227
rect 36 148 52 219
rect 90 194 123 202
rect 90 177 98 194
rect 115 177 123 194
rect 90 169 123 177
rect 36 133 87 148
rect 72 115 87 133
rect 108 115 123 169
rect 72 52 87 65
rect 108 52 123 65
<< polycont >>
rect 27 227 44 244
rect 98 237 115 254
rect 98 177 115 194
<< locali >>
rect 0 470 213 480
rect 0 442 28 470
rect 185 442 213 470
rect 0 432 213 442
rect 36 407 69 432
rect 36 323 44 407
rect 61 323 69 407
rect 36 315 69 323
rect 144 407 177 415
rect 144 323 152 407
rect 169 323 177 407
rect 90 254 123 262
rect 19 244 52 252
rect 19 227 27 244
rect 44 227 52 244
rect 90 237 98 254
rect 115 237 123 254
rect 90 229 123 237
rect 19 219 52 227
rect 90 194 123 202
rect 90 177 98 194
rect 115 177 123 194
rect 90 169 123 177
rect 144 115 177 323
rect 36 107 69 115
rect 36 73 44 107
rect 61 73 69 107
rect 36 48 69 73
rect 126 107 177 115
rect 126 73 134 107
rect 151 73 177 107
rect 126 65 177 73
rect 0 38 213 48
rect 0 10 12 38
rect 201 10 213 38
rect 0 0 213 10
<< labels >>
flabel ndiff 72 90 72 90 1 FreeSerif 8 0 0 0 S$
flabel pdiff 72 365 72 365 1 FreeSerif 8 0 0 0 S$
flabel ndiff 108 90 108 90 1 FreeSerif 8 0 0 0 S$
flabel locali 0 432 213 480 0 FreeSerif 80 0 0 0 VDD!
port 2 nsew
flabel locali 145 65 177 290 0 FreeSerif 80 0 0 0 Y
port 5 nsew
flabel locali 0 0 213 48 0 FreeSerif 80 0 0 0 GND!
port 3 nsew
flabel locali 19 219 52 252 0 FreeSerif 80 0 0 0 A
port 4 nsew
flabel locali 90 169 123 202 0 FreeSerif 80 0 0 0 EN
port 8 nsew
flabel locali 90 229 123 262 0 FreeSerif 80 0 0 0 ~EN
port 9 nsew
flabel pdiff 126 365 126 365 1 FreeSerif 8 0 0 0 S$
<< end >>
