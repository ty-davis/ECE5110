magic
tech sky130A
timestamp 1740425971
<< nwell >>
rect -2 197 323 488
<< nmos >>
rect 72 87 87 137
rect 126 87 141 137
rect 180 99 195 149
rect 234 99 249 149
<< pmos >>
rect 72 280 87 380
rect 126 280 141 380
rect 180 280 195 380
rect 234 280 249 380
<< ndiff >>
rect 155 137 180 149
rect 36 129 72 137
rect 36 95 44 129
rect 61 95 72 129
rect 36 87 72 95
rect 87 129 126 137
rect 87 95 98 129
rect 115 95 126 129
rect 87 87 126 95
rect 141 133 180 137
rect 141 99 151 133
rect 168 99 180 133
rect 195 141 234 149
rect 195 107 206 141
rect 223 107 234 141
rect 195 99 234 107
rect 249 141 285 149
rect 249 107 260 141
rect 277 107 285 141
rect 249 99 285 107
rect 141 87 172 99
<< pdiff >>
rect 36 372 72 380
rect 36 288 44 372
rect 61 288 72 372
rect 36 280 72 288
rect 87 372 126 380
rect 87 288 98 372
rect 115 288 126 372
rect 87 280 126 288
rect 141 372 180 380
rect 141 288 152 372
rect 169 288 180 372
rect 141 280 180 288
rect 195 372 234 380
rect 195 288 206 372
rect 223 288 234 372
rect 195 280 234 288
rect 249 372 285 380
rect 249 288 260 372
rect 277 288 285 372
rect 249 280 285 288
<< ndiffc >>
rect 44 95 61 129
rect 98 95 115 129
rect 151 99 168 133
rect 206 107 223 141
rect 260 107 277 141
<< pdiffc >>
rect 44 288 61 372
rect 98 288 115 372
rect 152 288 169 372
rect 206 288 223 372
rect 260 288 277 372
<< psubdiff >>
rect 0 10 12 38
rect 309 10 321 38
<< nsubdiff >>
rect 16 442 28 470
rect 293 442 305 470
<< psubdiffcont >>
rect 12 10 309 38
<< nsubdiffcont >>
rect 28 442 293 470
<< poly >>
rect 72 380 87 393
rect 126 380 141 393
rect 180 380 195 393
rect 234 380 249 393
rect 72 233 87 280
rect 54 225 87 233
rect 126 229 141 280
rect 180 229 195 280
rect 54 208 62 225
rect 79 208 87 225
rect 54 200 87 208
rect 72 137 87 200
rect 108 221 141 229
rect 108 204 116 221
rect 133 204 141 221
rect 108 196 141 204
rect 162 221 195 229
rect 162 204 170 221
rect 187 204 195 221
rect 162 196 195 204
rect 126 137 141 196
rect 180 149 195 196
rect 234 263 249 280
rect 234 255 282 263
rect 234 238 257 255
rect 274 238 282 255
rect 234 230 282 238
rect 234 149 249 230
rect 72 74 87 87
rect 126 74 141 87
rect 180 86 195 99
rect 234 86 249 99
<< polycont >>
rect 62 208 79 225
rect 116 204 133 221
rect 170 204 187 221
rect 257 238 274 255
<< locali >>
rect 0 470 321 480
rect 0 442 28 470
rect 293 442 321 470
rect 0 432 321 442
rect 36 372 69 432
rect 36 288 44 372
rect 61 288 69 372
rect 36 280 69 288
rect 90 398 231 415
rect 90 372 123 398
rect 90 288 98 372
rect 115 288 123 372
rect 90 280 123 288
rect 144 372 177 380
rect 144 288 152 372
rect 169 288 177 372
rect 144 263 177 288
rect 198 372 231 398
rect 198 288 206 372
rect 223 288 231 372
rect 198 280 231 288
rect 252 372 285 432
rect 252 288 260 372
rect 277 288 285 372
rect 252 280 285 288
rect 144 246 231 263
rect 54 225 87 233
rect 54 208 62 225
rect 79 208 87 225
rect 54 200 87 208
rect 108 221 141 229
rect 108 204 116 221
rect 133 204 141 221
rect 108 196 141 204
rect 162 221 195 229
rect 162 204 170 221
rect 187 204 195 221
rect 162 196 195 204
rect 212 202 231 246
rect 249 255 282 263
rect 249 238 257 255
rect 274 238 282 255
rect 249 230 282 238
rect 284 202 317 213
rect 212 180 317 202
rect 36 154 177 171
rect 212 168 231 180
rect 36 129 69 154
rect 36 95 44 129
rect 61 95 69 129
rect 36 87 69 95
rect 90 129 123 137
rect 90 95 98 129
rect 115 95 123 129
rect 90 48 123 95
rect 144 133 177 154
rect 144 99 151 133
rect 168 99 177 133
rect 198 141 231 168
rect 198 107 206 141
rect 223 107 231 141
rect 198 99 231 107
rect 252 141 285 149
rect 252 107 260 141
rect 277 107 285 141
rect 144 82 177 99
rect 252 82 285 107
rect 144 65 285 82
rect 0 38 321 48
rect 0 10 12 38
rect 309 10 321 38
rect 0 0 321 10
<< labels >>
flabel locali 0 0 321 48 0 FreeSerif 80 0 0 0 GND!
port 3 nsew
flabel locali 0 432 321 480 0 FreeSerif 80 0 0 0 VDD!
port 2 nsew
flabel pdiff 126 328 126 328 1 FreeSerif 8 0 0 0 S$
flabel pdiff 249 330 249 330 1 FreeSerif 8 0 0 0 S$
flabel pdiff 195 330 195 330 1 FreeSerif 8 0 0 0 S$
flabel pdiff 72 330 72 330 1 FreeSerif 8 0 0 0 S$
flabel ndiff 249 124 249 124 1 FreeSerif 8 0 0 0 S$
flabel ndiff 180 123 180 123 1 FreeSerif 8 0 0 0 S$
flabel locali 284 198 317 213 0 FreeSerif 80 0 0 0 Y
port 4 nsew
flabel ndiff 126 111 126 111 1 FreeSerif 8 0 0 0 S$
flabel ndiff 87 109 87 109 1 FreeSerif 8 0 0 0 S$
flabel locali 54 200 87 233 0 FreeSerif 80 0 0 0 C
port 11 nsew
flabel locali 108 196 141 229 0 FreeSerif 80 0 0 0 A
port 12 nsew
flabel locali 162 196 195 229 0 FreeSerif 80 0 0 0 B
port 14 nsew
flabel locali 249 230 282 263 0 FreeSerif 80 0 0 0 D
port 13 nsew
<< end >>
