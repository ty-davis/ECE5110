magic
tech sky130A
timestamp 1741762535
<< nwell >>
rect -2 197 856 488
<< nmos >>
rect 72 65 87 115
rect 126 65 141 115
rect 247 65 262 115
rect 361 65 376 115
rect 498 65 513 115
rect 552 65 567 115
rect 673 65 688 115
rect 787 65 802 115
<< pmos >>
rect 72 315 87 415
rect 126 315 141 415
rect 247 315 262 415
rect 361 315 376 415
rect 498 315 513 415
rect 552 315 567 415
rect 673 315 688 415
rect 787 315 802 415
<< ndiff >>
rect 36 107 72 115
rect 36 73 44 107
rect 61 73 72 107
rect 36 65 72 73
rect 87 107 126 115
rect 87 73 98 107
rect 115 73 126 107
rect 87 65 126 73
rect 141 107 177 115
rect 141 73 152 107
rect 169 73 177 107
rect 141 65 177 73
rect 211 107 247 115
rect 211 73 219 107
rect 236 73 247 107
rect 211 65 247 73
rect 262 107 298 115
rect 262 73 273 107
rect 290 73 298 107
rect 262 65 298 73
rect 325 107 361 115
rect 325 73 333 107
rect 350 73 361 107
rect 325 65 361 73
rect 376 107 412 115
rect 376 73 387 107
rect 404 73 412 107
rect 376 65 412 73
rect 462 107 498 115
rect 462 73 470 107
rect 487 73 498 107
rect 462 65 498 73
rect 513 107 552 115
rect 513 73 524 107
rect 541 73 552 107
rect 513 65 552 73
rect 567 107 603 115
rect 567 73 578 107
rect 595 73 603 107
rect 567 65 603 73
rect 637 107 673 115
rect 637 73 645 107
rect 662 73 673 107
rect 637 65 673 73
rect 688 107 724 115
rect 688 73 699 107
rect 716 73 724 107
rect 688 65 724 73
rect 751 107 787 115
rect 751 73 759 107
rect 776 73 787 107
rect 751 65 787 73
rect 802 107 838 115
rect 802 73 813 107
rect 830 73 838 107
rect 802 65 838 73
<< pdiff >>
rect 36 407 72 415
rect 36 323 44 407
rect 61 323 72 407
rect 36 315 72 323
rect 87 407 126 415
rect 87 323 98 407
rect 115 323 126 407
rect 87 315 126 323
rect 141 407 177 415
rect 141 323 152 407
rect 169 323 177 407
rect 141 315 177 323
rect 211 407 247 415
rect 211 323 219 407
rect 236 323 247 407
rect 211 315 247 323
rect 262 407 298 415
rect 262 323 273 407
rect 290 323 298 407
rect 262 315 298 323
rect 325 407 361 415
rect 325 323 333 407
rect 350 323 361 407
rect 325 315 361 323
rect 376 407 412 415
rect 376 323 387 407
rect 404 323 412 407
rect 376 315 412 323
rect 462 407 498 415
rect 462 323 470 407
rect 487 323 498 407
rect 462 315 498 323
rect 513 407 552 415
rect 513 323 524 407
rect 541 323 552 407
rect 513 315 552 323
rect 567 407 603 415
rect 567 323 578 407
rect 595 323 603 407
rect 567 315 603 323
rect 637 407 673 415
rect 637 323 645 407
rect 662 323 673 407
rect 637 315 673 323
rect 688 407 724 415
rect 688 323 699 407
rect 716 323 724 407
rect 688 315 724 323
rect 751 407 787 415
rect 751 323 759 407
rect 776 323 787 407
rect 751 315 787 323
rect 802 407 838 415
rect 802 323 813 407
rect 830 323 838 407
rect 802 315 838 323
<< ndiffc >>
rect 44 73 61 107
rect 98 73 115 107
rect 152 73 169 107
rect 219 73 236 107
rect 273 73 290 107
rect 333 73 350 107
rect 387 73 404 107
rect 470 73 487 107
rect 524 73 541 107
rect 578 73 595 107
rect 645 73 662 107
rect 699 73 716 107
rect 759 73 776 107
rect 813 73 830 107
<< pdiffc >>
rect 44 323 61 407
rect 98 323 115 407
rect 152 323 169 407
rect 219 323 236 407
rect 273 323 290 407
rect 333 323 350 407
rect 387 323 404 407
rect 470 323 487 407
rect 524 323 541 407
rect 578 323 595 407
rect 645 323 662 407
rect 699 323 716 407
rect 759 323 776 407
rect 813 323 830 407
<< psubdiff >>
rect 0 10 12 38
rect 842 10 854 38
<< nsubdiff >>
rect 16 442 28 470
rect 826 442 838 470
<< psubdiffcont >>
rect 12 10 842 38
<< nsubdiffcont >>
rect 28 442 826 470
<< poly >>
rect 72 415 87 428
rect 126 415 141 428
rect 247 415 262 428
rect 361 415 376 428
rect 498 415 513 428
rect 552 415 567 428
rect 673 415 688 428
rect 787 415 802 428
rect 72 224 87 315
rect 126 282 141 315
rect 126 274 159 282
rect 126 257 134 274
rect 151 257 159 274
rect 247 265 262 315
rect 126 249 159 257
rect 214 257 262 265
rect 361 261 376 315
rect 498 295 513 315
rect 480 287 513 295
rect 480 270 488 287
rect 505 270 513 287
rect 480 262 513 270
rect 214 240 222 257
rect 239 240 262 257
rect 214 232 262 240
rect 72 207 141 224
rect 115 199 141 207
rect 42 175 75 183
rect 42 158 50 175
rect 67 158 75 175
rect 126 182 141 199
rect 126 174 159 182
rect 42 150 87 158
rect 57 139 87 150
rect 72 115 87 139
rect 126 157 134 174
rect 151 157 159 174
rect 126 149 159 157
rect 126 115 141 149
rect 247 115 262 232
rect 328 253 376 261
rect 328 236 336 253
rect 353 236 376 253
rect 328 228 376 236
rect 552 228 567 315
rect 361 115 376 228
rect 483 213 567 228
rect 673 217 688 315
rect 787 261 802 315
rect 754 253 802 261
rect 754 236 762 253
rect 779 236 802 253
rect 754 228 802 236
rect 483 183 498 213
rect 640 209 688 217
rect 640 192 648 209
rect 665 192 688 209
rect 465 175 498 183
rect 465 158 473 175
rect 490 158 498 175
rect 465 150 498 158
rect 552 184 585 192
rect 640 184 688 192
rect 552 167 560 184
rect 577 167 585 184
rect 552 159 585 167
rect 478 135 513 150
rect 498 115 513 135
rect 552 115 567 159
rect 673 115 688 184
rect 787 115 802 228
rect 72 52 87 65
rect 126 52 141 65
rect 247 52 262 65
rect 361 52 376 65
rect 498 52 513 65
rect 552 52 567 65
rect 673 52 688 65
rect 787 52 802 65
<< polycont >>
rect 134 257 151 274
rect 488 270 505 287
rect 222 240 239 257
rect 50 158 67 175
rect 134 157 151 174
rect 336 236 353 253
rect 762 236 779 253
rect 648 192 665 209
rect 473 158 490 175
rect 560 167 577 184
<< locali >>
rect 0 470 854 480
rect 0 442 28 470
rect 826 442 854 470
rect 0 432 854 442
rect 36 407 69 415
rect 36 323 44 407
rect 61 323 69 407
rect 36 315 69 323
rect 90 407 123 415
rect 90 323 98 407
rect 115 323 123 407
rect 90 315 123 323
rect 144 407 177 415
rect 144 323 152 407
rect 169 323 177 407
rect 144 316 177 323
rect 211 407 244 432
rect 211 323 219 407
rect 236 323 244 407
rect 36 272 58 315
rect 20 256 58 272
rect 20 255 54 256
rect 7 247 40 255
rect 7 230 15 247
rect 32 230 40 247
rect 7 222 40 230
rect 90 232 107 315
rect 144 299 194 316
rect 211 315 244 323
rect 265 407 298 415
rect 265 323 273 407
rect 290 323 298 407
rect 126 274 159 282
rect 126 257 134 274
rect 151 257 159 274
rect 126 249 159 257
rect 90 224 128 232
rect 8 133 25 222
rect 90 207 103 224
rect 120 207 128 224
rect 92 199 128 207
rect 42 175 75 183
rect 42 158 50 175
rect 67 158 75 175
rect 42 150 75 158
rect 8 115 69 133
rect 92 119 109 199
rect 176 197 194 299
rect 214 257 247 265
rect 214 240 222 257
rect 239 240 247 257
rect 214 232 247 240
rect 265 251 298 323
rect 325 407 358 432
rect 325 323 333 407
rect 350 323 358 407
rect 325 315 358 323
rect 379 407 412 415
rect 379 323 387 407
rect 404 323 412 407
rect 462 407 495 415
rect 462 332 470 407
rect 328 253 361 261
rect 328 251 336 253
rect 265 236 336 251
rect 353 236 361 253
rect 265 228 361 236
rect 126 174 159 182
rect 126 157 134 174
rect 151 157 159 174
rect 126 149 159 157
rect 176 165 193 197
rect 176 157 209 165
rect 176 140 184 157
rect 201 140 209 157
rect 176 132 209 140
rect 36 107 69 115
rect 36 73 44 107
rect 61 73 69 107
rect 36 65 69 73
rect 90 107 123 119
rect 90 73 98 107
rect 115 73 123 107
rect 90 65 123 73
rect 144 115 194 132
rect 144 107 177 115
rect 144 73 152 107
rect 169 73 177 107
rect 144 65 177 73
rect 211 107 244 115
rect 211 73 219 107
rect 236 73 244 107
rect 211 48 244 73
rect 265 107 298 228
rect 379 157 412 323
rect 445 323 470 332
rect 487 323 495 407
rect 445 315 495 323
rect 516 407 549 415
rect 516 323 524 407
rect 541 323 549 407
rect 516 315 549 323
rect 445 255 462 315
rect 480 287 513 295
rect 480 270 488 287
rect 505 270 513 287
rect 480 262 513 270
rect 379 140 387 157
rect 404 140 412 157
rect 265 73 273 107
rect 290 73 298 107
rect 265 65 298 73
rect 325 107 358 115
rect 325 73 333 107
rect 350 73 358 107
rect 325 48 358 73
rect 379 107 412 140
rect 429 247 462 255
rect 429 230 437 247
rect 454 230 462 247
rect 532 261 549 315
rect 570 407 603 415
rect 570 323 578 407
rect 595 323 603 407
rect 570 316 603 323
rect 637 407 670 432
rect 637 323 645 407
rect 662 323 670 407
rect 570 299 620 316
rect 637 315 670 323
rect 691 407 724 415
rect 691 323 699 407
rect 716 323 724 407
rect 532 253 565 261
rect 532 245 540 253
rect 429 222 462 230
rect 516 236 540 245
rect 557 236 565 253
rect 516 228 565 236
rect 429 133 446 222
rect 465 175 498 183
rect 465 158 473 175
rect 490 158 498 175
rect 465 150 498 158
rect 429 115 495 133
rect 379 73 387 107
rect 404 73 412 107
rect 379 65 412 73
rect 462 107 495 115
rect 462 73 470 107
rect 487 73 495 107
rect 462 65 495 73
rect 516 115 533 228
rect 552 184 585 192
rect 552 167 560 184
rect 577 167 585 184
rect 552 159 585 167
rect 602 165 620 299
rect 691 251 724 323
rect 751 407 784 432
rect 751 323 759 407
rect 776 323 784 407
rect 751 315 784 323
rect 805 407 838 415
rect 805 323 813 407
rect 830 323 838 407
rect 754 253 787 261
rect 754 251 762 253
rect 691 236 762 251
rect 779 236 787 253
rect 691 228 787 236
rect 640 209 673 217
rect 640 192 648 209
rect 665 192 673 209
rect 640 184 673 192
rect 602 157 635 165
rect 602 140 610 157
rect 627 140 635 157
rect 602 132 635 140
rect 570 115 620 132
rect 691 115 708 228
rect 805 157 838 323
rect 805 140 813 157
rect 830 140 838 157
rect 516 107 549 115
rect 516 73 524 107
rect 541 73 549 107
rect 516 65 549 73
rect 570 107 603 115
rect 570 73 578 107
rect 595 73 603 107
rect 570 65 603 73
rect 637 107 670 115
rect 637 73 645 107
rect 662 73 670 107
rect 637 48 670 73
rect 691 107 724 115
rect 691 73 699 107
rect 716 73 724 107
rect 691 65 724 73
rect 751 107 784 115
rect 751 73 759 107
rect 776 73 784 107
rect 751 48 784 73
rect 805 107 838 140
rect 805 73 813 107
rect 830 73 838 107
rect 805 65 838 73
rect 0 38 854 48
rect 0 10 12 38
rect 842 10 854 38
rect 0 0 854 10
<< viali >>
rect 15 230 32 247
rect 134 257 151 274
rect 103 207 120 224
rect 50 158 67 175
rect 222 240 239 257
rect 336 236 353 253
rect 134 157 151 174
rect 184 140 201 157
rect 488 270 505 287
rect 387 140 404 157
rect 437 230 454 247
rect 540 236 557 253
rect 473 158 490 175
rect 560 167 577 184
rect 648 192 665 209
rect 610 140 627 157
rect 813 140 830 157
<< metal1 >>
rect 145 287 513 295
rect 145 282 488 287
rect 126 281 488 282
rect 126 274 159 281
rect 126 263 134 274
rect 54 257 134 263
rect 151 257 159 274
rect 480 270 488 281
rect 505 270 513 287
rect 7 247 40 255
rect 7 230 15 247
rect 32 230 40 247
rect 7 222 40 230
rect 54 249 159 257
rect 214 257 247 265
rect 480 262 513 270
rect 54 183 70 249
rect 214 240 222 257
rect 239 240 247 257
rect 214 232 247 240
rect 328 255 361 261
rect 328 253 462 255
rect 328 236 336 253
rect 353 247 462 253
rect 353 237 437 247
rect 353 236 361 237
rect 95 224 228 232
rect 328 228 361 236
rect 429 230 437 237
rect 454 230 462 247
rect 95 207 103 224
rect 120 216 228 224
rect 429 222 462 230
rect 120 207 128 216
rect 95 199 128 207
rect 499 211 513 262
rect 532 253 565 261
rect 532 236 540 253
rect 557 244 565 253
rect 557 236 640 244
rect 532 229 640 236
rect 532 228 565 229
rect 625 217 640 229
rect 499 197 552 211
rect 625 209 673 217
rect 625 201 648 209
rect 145 183 465 193
rect 538 192 552 197
rect 640 192 648 201
rect 665 192 673 209
rect 538 184 585 192
rect 640 184 673 192
rect 42 175 75 183
rect 145 182 498 183
rect 42 158 50 175
rect 67 158 75 175
rect 42 150 75 158
rect 126 179 498 182
rect 126 174 159 179
rect 126 157 134 174
rect 151 157 159 174
rect 451 175 498 179
rect 538 177 560 184
rect 451 167 473 175
rect 126 149 159 157
rect 176 157 412 165
rect 176 140 184 157
rect 201 150 387 157
rect 201 140 209 150
rect 176 132 209 140
rect 379 140 387 150
rect 404 140 412 157
rect 465 158 473 167
rect 490 158 498 175
rect 552 167 560 177
rect 577 167 585 184
rect 552 159 585 167
rect 465 150 498 158
rect 602 157 838 165
rect 379 132 412 140
rect 602 140 610 157
rect 627 150 813 157
rect 627 140 635 150
rect 728 149 773 150
rect 602 132 635 140
rect 805 140 813 150
rect 830 140 838 157
rect 805 132 838 140
<< labels >>
flabel pdiff 247 365 247 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 361 365 361 365 1 FreeSerif 8 0 0 0 S$
flabel ndiff 361 90 361 90 1 FreeSerif 8 0 0 0 S$
flabel pdiff 87 366 87 366 1 FreeSerif 8 0 0 0 S$
flabel pdiff 141 366 141 366 1 FreeSerif 8 0 0 0 S$
flabel ndiff 141 90 141 90 1 FreeSerif 8 0 0 0 S$
flabel ndiff 87 90 87 90 1 FreeSerif 8 0 0 0 S$
flabel ndiff 247 90 247 90 1 FreeSerif 8 0 0 0 S$
flabel pdiff 673 365 673 365 1 FreeSerif 8 0 0 0 S$
flabel ndiff 673 90 673 90 1 FreeSerif 8 0 0 0 S$
flabel pdiff 787 365 787 365 1 FreeSerif 8 0 0 0 S$
flabel ndiff 787 90 787 90 1 FreeSerif 8 0 0 0 S$
flabel pdiff 513 366 513 366 1 FreeSerif 8 0 0 0 S$
flabel pdiff 567 366 567 366 1 FreeSerif 8 0 0 0 S$
flabel ndiff 567 90 567 90 1 FreeSerif 8 0 0 0 S$
flabel ndiff 513 90 513 90 1 FreeSerif 8 0 0 0 S$
flabel locali 0 432 854 480 0 FreeSerif 80 0 0 0 VDD!
port 15 nsew
flabel locali 126 149 134 182 0 FreeSerif 80 0 0 0 CLK
port 2 nsew
flabel locali 7 222 40 255 0 FreeSerif 80 0 0 0 D
port 0 nsew
flabel locali 0 0 854 48 0 FreeSerif 80 0 0 0 GND!
port 16 nsew
flabel locali 126 249 134 282 0 FreeSerif 80 0 0 0 ~CLK
port 1 nsew
flabel locali 805 182 838 219 0 FreeSerif 80 0 0 0 ~Q
port 3 nsew
flabel locali 754 228 787 261 0 FreeSerif 80 0 0 0 Q
port 4 nsew
<< end >>
