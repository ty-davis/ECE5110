magic
tech sky130A
magscale 1 2
timestamp 1745353766
<< error_p >>
rect 242 -222 247 -136
<< nwell >>
rect -36 -492 1880 254
<< nmos >>
rect 258 352 292 438
rect 490 352 524 438
rect 722 352 756 438
rect 954 352 988 438
rect 1186 352 1220 438
rect 1418 352 1452 438
rect 1650 352 1684 438
<< pmos >>
rect 258 132 292 218
rect 490 132 524 218
rect 722 132 756 218
rect 954 132 988 218
rect 1186 132 1220 218
rect 1418 132 1452 218
rect 1650 132 1684 218
rect 314 -222 348 -136
rect 434 -222 468 -136
rect 546 -222 580 -136
rect 666 -222 700 -136
rect 778 -222 812 -136
rect 898 -222 932 -136
rect 1010 -222 1044 -136
rect 1130 -222 1164 -136
rect 1242 -222 1276 -136
rect 1362 -222 1396 -136
rect 1474 -222 1508 -136
rect 1594 -222 1628 -136
rect 1706 -222 1740 -136
rect 202 -362 236 -276
rect 314 -362 348 -276
rect 434 -362 468 -276
rect 546 -362 580 -276
rect 666 -362 700 -276
rect 778 -362 812 -276
rect 898 -362 932 -276
rect 1010 -362 1044 -276
rect 1130 -362 1164 -276
rect 1242 -362 1276 -276
rect 1362 -362 1396 -276
rect 1474 -362 1508 -276
rect 1594 -362 1628 -276
rect 1706 -362 1740 -276
<< ndiff >>
rect 186 422 258 438
rect 186 368 202 422
rect 236 368 258 422
rect 186 352 258 368
rect 292 422 364 438
rect 292 368 314 422
rect 348 368 364 422
rect 292 352 364 368
rect 418 422 490 438
rect 418 368 434 422
rect 468 368 490 422
rect 418 352 490 368
rect 524 422 596 438
rect 524 368 546 422
rect 580 368 596 422
rect 524 352 596 368
rect 650 422 722 438
rect 650 368 666 422
rect 700 368 722 422
rect 650 352 722 368
rect 756 422 828 438
rect 756 368 778 422
rect 812 368 828 422
rect 756 352 828 368
rect 882 422 954 438
rect 882 368 898 422
rect 932 368 954 422
rect 882 352 954 368
rect 988 422 1060 438
rect 988 368 1010 422
rect 1044 368 1060 422
rect 988 352 1060 368
rect 1114 422 1186 438
rect 1114 368 1130 422
rect 1164 368 1186 422
rect 1114 352 1186 368
rect 1220 422 1292 438
rect 1220 368 1242 422
rect 1276 368 1292 422
rect 1220 352 1292 368
rect 1346 422 1418 438
rect 1346 368 1362 422
rect 1396 368 1418 422
rect 1346 352 1418 368
rect 1452 422 1524 438
rect 1452 368 1474 422
rect 1508 368 1524 422
rect 1452 352 1524 368
rect 1578 422 1650 438
rect 1578 368 1594 422
rect 1628 368 1650 422
rect 1578 352 1650 368
rect 1684 422 1756 438
rect 1684 368 1706 422
rect 1740 368 1756 422
rect 1684 352 1756 368
<< pdiff >>
rect 186 202 258 218
rect 186 148 202 202
rect 236 148 258 202
rect 186 132 258 148
rect 292 202 364 218
rect 292 148 314 202
rect 348 148 364 202
rect 292 132 364 148
rect 418 202 490 218
rect 418 148 434 202
rect 468 148 490 202
rect 418 132 490 148
rect 524 202 596 218
rect 524 148 546 202
rect 580 148 596 202
rect 524 132 596 148
rect 650 202 722 218
rect 650 148 666 202
rect 700 148 722 202
rect 650 132 722 148
rect 756 202 828 218
rect 756 148 778 202
rect 812 148 828 202
rect 756 132 828 148
rect 882 202 954 218
rect 882 148 898 202
rect 932 148 954 202
rect 882 132 954 148
rect 988 202 1060 218
rect 988 148 1010 202
rect 1044 148 1060 202
rect 988 132 1060 148
rect 1114 202 1186 218
rect 1114 148 1130 202
rect 1164 148 1186 202
rect 1114 132 1186 148
rect 1220 202 1292 218
rect 1220 148 1242 202
rect 1276 148 1292 202
rect 1220 132 1292 148
rect 1346 202 1418 218
rect 1346 148 1362 202
rect 1396 148 1418 202
rect 1346 132 1418 148
rect 1452 202 1524 218
rect 1452 148 1474 202
rect 1508 148 1524 202
rect 1452 132 1524 148
rect 1578 202 1650 218
rect 1578 148 1594 202
rect 1628 148 1650 202
rect 1578 132 1650 148
rect 1684 202 1756 218
rect 1684 148 1706 202
rect 1740 148 1756 202
rect 1684 132 1756 148
rect 242 -152 314 -136
rect 242 -206 258 -152
rect 292 -206 314 -152
rect 242 -222 314 -206
rect 348 -152 434 -136
rect 348 -206 370 -152
rect 412 -206 434 -152
rect 348 -222 434 -206
rect 468 -152 546 -136
rect 468 -206 490 -152
rect 524 -206 546 -152
rect 468 -222 546 -206
rect 580 -152 666 -136
rect 580 -206 602 -152
rect 644 -206 666 -152
rect 580 -222 666 -206
rect 700 -152 778 -136
rect 700 -206 722 -152
rect 756 -206 778 -152
rect 700 -222 778 -206
rect 812 -152 898 -136
rect 812 -206 834 -152
rect 876 -206 898 -152
rect 812 -222 898 -206
rect 932 -152 1010 -136
rect 932 -206 954 -152
rect 988 -206 1010 -152
rect 932 -222 1010 -206
rect 1044 -152 1130 -136
rect 1044 -206 1066 -152
rect 1108 -206 1130 -152
rect 1044 -222 1130 -206
rect 1164 -152 1242 -136
rect 1164 -206 1186 -152
rect 1220 -206 1242 -152
rect 1164 -222 1242 -206
rect 1276 -152 1362 -136
rect 1276 -206 1298 -152
rect 1340 -206 1362 -152
rect 1276 -222 1362 -206
rect 1396 -152 1474 -136
rect 1396 -206 1418 -152
rect 1452 -206 1474 -152
rect 1396 -222 1474 -206
rect 1508 -152 1594 -136
rect 1508 -206 1530 -152
rect 1572 -206 1594 -152
rect 1508 -222 1594 -206
rect 1628 -152 1706 -136
rect 1628 -206 1650 -152
rect 1684 -206 1706 -152
rect 1628 -222 1706 -206
rect 1740 -152 1820 -136
rect 1740 -206 1762 -152
rect 1804 -206 1820 -152
rect 1740 -222 1820 -206
rect 130 -292 202 -276
rect 130 -346 146 -292
rect 180 -346 202 -292
rect 130 -362 202 -346
rect 236 -292 314 -276
rect 236 -346 258 -292
rect 292 -346 314 -292
rect 236 -362 314 -346
rect 348 -292 434 -276
rect 348 -346 370 -292
rect 412 -346 434 -292
rect 348 -362 434 -346
rect 468 -292 546 -276
rect 468 -346 490 -292
rect 524 -346 546 -292
rect 468 -362 546 -346
rect 580 -292 666 -276
rect 580 -346 602 -292
rect 644 -346 666 -292
rect 580 -362 666 -346
rect 700 -292 778 -276
rect 700 -346 722 -292
rect 756 -346 778 -292
rect 700 -362 778 -346
rect 812 -292 898 -276
rect 812 -346 834 -292
rect 876 -346 898 -292
rect 812 -362 898 -346
rect 932 -292 1010 -276
rect 932 -346 954 -292
rect 988 -346 1010 -292
rect 932 -362 1010 -346
rect 1044 -292 1130 -276
rect 1044 -346 1066 -292
rect 1108 -346 1130 -292
rect 1044 -362 1130 -346
rect 1164 -292 1242 -276
rect 1164 -346 1186 -292
rect 1220 -346 1242 -292
rect 1164 -362 1242 -346
rect 1276 -292 1362 -276
rect 1276 -346 1298 -292
rect 1340 -346 1362 -292
rect 1276 -362 1362 -346
rect 1396 -292 1474 -276
rect 1396 -346 1418 -292
rect 1452 -346 1474 -292
rect 1396 -362 1474 -346
rect 1508 -292 1594 -276
rect 1508 -346 1530 -292
rect 1572 -346 1594 -292
rect 1508 -362 1594 -346
rect 1628 -292 1706 -276
rect 1628 -346 1650 -292
rect 1684 -346 1706 -292
rect 1628 -362 1706 -346
rect 1740 -292 1820 -276
rect 1740 -346 1762 -292
rect 1804 -346 1820 -292
rect 1740 -362 1820 -346
<< ndiffc >>
rect 202 368 236 422
rect 314 368 348 422
rect 434 368 468 422
rect 546 368 580 422
rect 666 368 700 422
rect 778 368 812 422
rect 898 368 932 422
rect 1010 368 1044 422
rect 1130 368 1164 422
rect 1242 368 1276 422
rect 1362 368 1396 422
rect 1474 368 1508 422
rect 1594 368 1628 422
rect 1706 368 1740 422
<< pdiffc >>
rect 202 148 236 202
rect 314 148 348 202
rect 434 148 468 202
rect 546 148 580 202
rect 666 148 700 202
rect 778 148 812 202
rect 898 148 932 202
rect 1010 148 1044 202
rect 1130 148 1164 202
rect 1242 148 1276 202
rect 1362 148 1396 202
rect 1474 148 1508 202
rect 1594 148 1628 202
rect 1706 148 1740 202
rect 258 -206 292 -152
rect 370 -206 412 -152
rect 490 -206 524 -152
rect 602 -206 644 -152
rect 722 -206 756 -152
rect 834 -206 876 -152
rect 954 -206 988 -152
rect 1066 -206 1108 -152
rect 1186 -206 1220 -152
rect 1298 -206 1340 -152
rect 1418 -206 1452 -152
rect 1530 -206 1572 -152
rect 1650 -206 1684 -152
rect 1762 -206 1804 -152
rect 146 -346 180 -292
rect 258 -346 292 -292
rect 370 -346 412 -292
rect 490 -346 524 -292
rect 602 -346 644 -292
rect 722 -346 756 -292
rect 834 -346 876 -292
rect 954 -346 988 -292
rect 1066 -346 1108 -292
rect 1186 -346 1220 -292
rect 1298 -346 1340 -292
rect 1418 -346 1452 -292
rect 1530 -346 1572 -292
rect 1650 -346 1684 -292
rect 1762 -346 1804 -292
<< psubdiff >>
rect 24 492 48 548
rect 1820 492 1844 548
<< nsubdiff >>
rect 24 22 48 78
rect 1820 22 1844 78
rect 20 -56 76 -32
rect 20 -426 22 -56
rect 20 -450 76 -426
<< psubdiffcont >>
rect 48 492 1820 548
<< nsubdiffcont >>
rect 48 22 1820 78
rect 22 -426 76 -56
<< poly >>
rect 258 438 292 464
rect 490 438 524 464
rect 722 438 756 464
rect 954 438 988 464
rect 1186 438 1220 464
rect 1418 438 1452 464
rect 1650 438 1684 464
rect 258 318 292 352
rect 490 318 524 352
rect 722 318 756 352
rect 954 318 988 352
rect 1186 318 1220 352
rect 1418 318 1452 352
rect 1650 318 1684 352
rect 258 302 364 318
rect 258 268 314 302
rect 348 268 364 302
rect 258 252 364 268
rect 490 302 596 318
rect 490 268 546 302
rect 580 268 596 302
rect 490 252 596 268
rect 722 302 828 318
rect 722 268 778 302
rect 812 268 828 302
rect 722 252 828 268
rect 954 302 1060 318
rect 954 268 1010 302
rect 1044 268 1060 302
rect 954 252 1060 268
rect 1186 302 1292 318
rect 1186 268 1242 302
rect 1276 268 1292 302
rect 1186 252 1292 268
rect 1418 302 1524 318
rect 1418 268 1474 302
rect 1508 268 1524 302
rect 1418 252 1524 268
rect 1650 302 1756 318
rect 1650 268 1706 302
rect 1740 268 1756 302
rect 1650 252 1756 268
rect 258 218 292 252
rect 490 218 524 252
rect 722 218 756 252
rect 954 218 988 252
rect 1186 218 1220 252
rect 1418 218 1452 252
rect 1650 218 1684 252
rect 258 106 292 132
rect 490 106 524 132
rect 722 106 756 132
rect 954 106 988 132
rect 1186 106 1220 132
rect 1418 106 1452 132
rect 1650 106 1684 132
rect 186 -48 252 -32
rect 186 -82 202 -48
rect 236 -82 252 -48
rect 186 -98 252 -82
rect 298 -48 364 -32
rect 298 -82 314 -48
rect 348 -82 364 -48
rect 298 -98 364 -82
rect 418 -48 484 -32
rect 418 -82 434 -48
rect 468 -82 484 -48
rect 418 -98 484 -82
rect 530 -48 596 -32
rect 530 -82 546 -48
rect 580 -82 596 -48
rect 530 -98 596 -82
rect 650 -48 716 -32
rect 650 -82 666 -48
rect 700 -82 716 -48
rect 650 -98 716 -82
rect 762 -48 828 -32
rect 762 -82 778 -48
rect 812 -82 828 -48
rect 762 -98 828 -82
rect 882 -48 948 -32
rect 882 -82 898 -48
rect 932 -82 948 -48
rect 882 -98 948 -82
rect 994 -48 1060 -32
rect 994 -82 1010 -48
rect 1044 -82 1060 -48
rect 994 -98 1060 -82
rect 1114 -48 1180 -32
rect 1114 -82 1130 -48
rect 1164 -82 1180 -48
rect 1114 -98 1180 -82
rect 1226 -48 1292 -32
rect 1226 -82 1242 -48
rect 1276 -82 1292 -48
rect 1226 -98 1292 -82
rect 1346 -48 1412 -32
rect 1346 -82 1362 -48
rect 1396 -82 1412 -48
rect 1346 -98 1412 -82
rect 1458 -48 1524 -32
rect 1458 -82 1474 -48
rect 1508 -82 1524 -48
rect 1458 -98 1524 -82
rect 1578 -48 1644 -32
rect 1578 -82 1594 -48
rect 1628 -82 1644 -48
rect 1578 -98 1644 -82
rect 1690 -48 1756 -32
rect 1690 -82 1706 -48
rect 1740 -82 1756 -48
rect 1690 -98 1756 -82
rect 202 -114 236 -98
rect 202 -238 232 -114
rect 314 -136 348 -98
rect 434 -136 468 -98
rect 546 -136 580 -98
rect 666 -136 700 -98
rect 778 -136 812 -98
rect 898 -136 932 -98
rect 1010 -136 1044 -98
rect 1130 -136 1164 -98
rect 1242 -136 1276 -98
rect 1362 -136 1396 -98
rect 1474 -136 1508 -98
rect 1594 -136 1628 -98
rect 1706 -136 1740 -98
rect 202 -276 236 -238
rect 314 -276 348 -222
rect 434 -276 468 -222
rect 546 -276 580 -222
rect 666 -276 700 -222
rect 778 -276 812 -222
rect 898 -276 932 -222
rect 1010 -276 1044 -222
rect 1130 -276 1164 -222
rect 1242 -276 1276 -222
rect 1362 -276 1396 -222
rect 1474 -276 1508 -222
rect 1594 -276 1628 -222
rect 1706 -276 1740 -222
rect 202 -388 236 -362
rect 314 -388 348 -362
rect 434 -388 468 -362
rect 546 -388 580 -362
rect 666 -388 700 -362
rect 778 -388 812 -362
rect 898 -388 932 -362
rect 1010 -388 1044 -362
rect 1130 -388 1164 -362
rect 1242 -388 1276 -362
rect 1362 -388 1396 -362
rect 1474 -388 1508 -362
rect 1594 -388 1628 -362
rect 1706 -388 1740 -362
<< polycont >>
rect 314 268 348 302
rect 546 268 580 302
rect 778 268 812 302
rect 1010 268 1044 302
rect 1242 268 1276 302
rect 1474 268 1508 302
rect 1706 268 1740 302
rect 202 -82 236 -48
rect 314 -82 348 -48
rect 434 -82 468 -48
rect 546 -82 580 -48
rect 666 -82 700 -48
rect 778 -82 812 -48
rect 898 -82 932 -48
rect 1010 -82 1044 -48
rect 1130 -82 1164 -48
rect 1242 -82 1276 -48
rect 1362 -82 1396 -48
rect 1474 -82 1508 -48
rect 1594 -82 1628 -48
rect 1706 -82 1740 -48
<< locali >>
rect 0 548 1876 568
rect 0 492 48 548
rect 1820 492 1876 548
rect 0 472 1876 492
rect 186 422 252 438
rect 186 368 202 422
rect 236 368 252 422
rect 186 202 252 368
rect 298 422 364 472
rect 298 368 314 422
rect 348 368 364 422
rect 298 352 364 368
rect 418 422 484 438
rect 418 368 434 422
rect 468 368 484 422
rect 292 302 364 318
rect 292 268 314 302
rect 348 268 364 302
rect 292 252 364 268
rect 186 148 202 202
rect 236 148 252 202
rect 186 132 252 148
rect 298 202 364 218
rect 298 148 314 202
rect 348 148 364 202
rect 298 98 364 148
rect 418 202 484 368
rect 530 422 596 472
rect 530 368 546 422
rect 580 368 596 422
rect 530 352 596 368
rect 650 422 716 438
rect 650 368 666 422
rect 700 368 716 422
rect 524 302 596 318
rect 524 268 546 302
rect 580 268 596 302
rect 524 252 596 268
rect 418 148 434 202
rect 468 148 484 202
rect 418 132 484 148
rect 530 202 596 218
rect 530 148 546 202
rect 580 148 596 202
rect 530 98 596 148
rect 650 202 716 368
rect 762 422 828 472
rect 762 368 778 422
rect 812 368 828 422
rect 762 352 828 368
rect 882 422 948 438
rect 882 368 898 422
rect 932 368 948 422
rect 756 302 828 318
rect 756 268 778 302
rect 812 268 828 302
rect 756 252 828 268
rect 650 148 666 202
rect 700 148 716 202
rect 650 132 716 148
rect 762 202 828 218
rect 762 148 778 202
rect 812 148 828 202
rect 762 98 828 148
rect 882 202 948 368
rect 994 422 1060 472
rect 994 368 1010 422
rect 1044 368 1060 422
rect 994 352 1060 368
rect 1114 422 1180 438
rect 1114 368 1130 422
rect 1164 368 1180 422
rect 988 302 1060 318
rect 988 268 1010 302
rect 1044 268 1060 302
rect 988 252 1060 268
rect 882 148 898 202
rect 932 148 948 202
rect 882 132 948 148
rect 994 202 1060 218
rect 994 148 1010 202
rect 1044 148 1060 202
rect 994 98 1060 148
rect 1114 202 1180 368
rect 1226 422 1292 472
rect 1226 368 1242 422
rect 1276 368 1292 422
rect 1226 352 1292 368
rect 1346 422 1412 438
rect 1346 368 1362 422
rect 1396 368 1412 422
rect 1220 302 1292 318
rect 1220 268 1242 302
rect 1276 268 1292 302
rect 1220 252 1292 268
rect 1114 148 1130 202
rect 1164 148 1180 202
rect 1114 132 1180 148
rect 1226 202 1292 218
rect 1226 148 1242 202
rect 1276 148 1292 202
rect 1226 98 1292 148
rect 1346 202 1412 368
rect 1458 422 1524 472
rect 1458 368 1474 422
rect 1508 368 1524 422
rect 1458 352 1524 368
rect 1578 422 1644 438
rect 1578 368 1594 422
rect 1628 368 1644 422
rect 1452 302 1524 318
rect 1452 268 1474 302
rect 1508 268 1524 302
rect 1452 252 1524 268
rect 1346 148 1362 202
rect 1396 148 1412 202
rect 1346 132 1412 148
rect 1458 202 1524 218
rect 1458 148 1474 202
rect 1508 148 1524 202
rect 1458 98 1524 148
rect 1578 202 1644 368
rect 1690 422 1756 472
rect 1690 368 1706 422
rect 1740 368 1756 422
rect 1690 352 1756 368
rect 1684 302 1756 318
rect 1684 268 1706 302
rect 1740 268 1756 302
rect 1684 252 1756 268
rect 1578 148 1594 202
rect 1628 148 1644 202
rect 1578 132 1644 148
rect 1690 202 1756 218
rect 1690 148 1706 202
rect 1740 148 1756 202
rect 1690 98 1756 148
rect 0 78 1876 98
rect 0 22 48 78
rect 1820 22 1876 78
rect 0 2 1876 22
rect 0 -56 96 2
rect 0 -426 22 -56
rect 76 -136 96 -56
rect 186 -48 252 -32
rect 186 -82 202 -48
rect 236 -82 252 -48
rect 186 -98 252 -82
rect 298 -48 364 -32
rect 298 -82 314 -48
rect 348 -82 364 -48
rect 298 -98 364 -82
rect 418 -48 484 -32
rect 418 -82 434 -48
rect 468 -82 484 -48
rect 418 -98 484 -82
rect 530 -48 596 -32
rect 530 -82 546 -48
rect 580 -82 596 -48
rect 530 -98 596 -82
rect 650 -48 716 -32
rect 650 -82 666 -48
rect 700 -82 716 -48
rect 650 -98 716 -82
rect 762 -48 828 -32
rect 762 -82 778 -48
rect 812 -82 828 -48
rect 762 -98 828 -82
rect 882 -48 948 -32
rect 882 -82 898 -48
rect 932 -82 948 -48
rect 882 -98 948 -82
rect 994 -48 1060 -32
rect 994 -82 1010 -48
rect 1044 -82 1060 -48
rect 994 -98 1060 -82
rect 1114 -48 1180 -32
rect 1114 -82 1130 -48
rect 1164 -82 1180 -48
rect 1114 -98 1180 -82
rect 1226 -48 1292 -32
rect 1226 -82 1242 -48
rect 1276 -82 1292 -48
rect 1226 -98 1292 -82
rect 1346 -48 1412 -32
rect 1346 -82 1362 -48
rect 1396 -82 1412 -48
rect 1346 -98 1412 -82
rect 1458 -48 1524 -32
rect 1458 -82 1474 -48
rect 1508 -82 1524 -48
rect 1458 -98 1524 -82
rect 1578 -48 1644 -32
rect 1578 -82 1594 -48
rect 1628 -82 1644 -48
rect 1578 -98 1644 -82
rect 1690 -48 1756 -32
rect 1690 -82 1706 -48
rect 1740 -82 1756 -48
rect 1690 -98 1756 -82
rect 76 -152 308 -136
rect 76 -206 258 -152
rect 292 -206 308 -152
rect 76 -222 308 -206
rect 354 -152 428 -136
rect 354 -206 370 -152
rect 412 -206 428 -152
rect 354 -222 428 -206
rect 474 -152 540 -136
rect 474 -206 490 -152
rect 524 -206 540 -152
rect 474 -222 540 -206
rect 586 -152 660 -136
rect 586 -206 602 -152
rect 644 -206 660 -152
rect 586 -222 660 -206
rect 706 -152 772 -136
rect 706 -206 722 -152
rect 756 -206 772 -152
rect 706 -222 772 -206
rect 818 -152 892 -136
rect 818 -206 834 -152
rect 876 -206 892 -152
rect 818 -222 892 -206
rect 938 -152 1004 -136
rect 938 -206 954 -152
rect 988 -206 1004 -152
rect 938 -222 1004 -206
rect 1050 -152 1124 -136
rect 1050 -206 1066 -152
rect 1108 -206 1124 -152
rect 1050 -222 1124 -206
rect 1170 -152 1236 -136
rect 1170 -206 1186 -152
rect 1220 -206 1236 -152
rect 1170 -222 1236 -206
rect 1282 -152 1356 -136
rect 1282 -206 1298 -152
rect 1340 -206 1356 -152
rect 1282 -222 1356 -206
rect 1402 -152 1468 -136
rect 1402 -206 1418 -152
rect 1452 -206 1468 -152
rect 1402 -222 1468 -206
rect 1514 -152 1588 -136
rect 1514 -206 1530 -152
rect 1572 -206 1588 -152
rect 1514 -222 1588 -206
rect 1634 -152 1700 -136
rect 1634 -206 1650 -152
rect 1684 -206 1700 -152
rect 1634 -222 1700 -206
rect 1746 -152 1820 -136
rect 1746 -206 1762 -152
rect 1804 -206 1820 -152
rect 1746 -222 1820 -206
rect 76 -276 96 -222
rect 76 -292 196 -276
rect 76 -346 146 -292
rect 180 -346 196 -292
rect 76 -362 196 -346
rect 242 -292 308 -276
rect 242 -346 258 -292
rect 292 -346 308 -292
rect 242 -362 308 -346
rect 354 -292 428 -276
rect 354 -346 370 -292
rect 412 -346 428 -292
rect 354 -362 428 -346
rect 474 -292 540 -276
rect 474 -346 490 -292
rect 524 -346 540 -292
rect 474 -362 540 -346
rect 586 -292 660 -276
rect 586 -346 602 -292
rect 644 -346 660 -292
rect 586 -362 660 -346
rect 706 -292 772 -276
rect 706 -346 722 -292
rect 756 -346 772 -292
rect 706 -362 772 -346
rect 818 -292 892 -276
rect 818 -346 834 -292
rect 876 -346 892 -292
rect 818 -362 892 -346
rect 938 -292 1004 -276
rect 938 -346 954 -292
rect 988 -346 1004 -292
rect 938 -362 1004 -346
rect 1050 -292 1124 -276
rect 1050 -346 1066 -292
rect 1108 -346 1124 -292
rect 1050 -362 1124 -346
rect 1170 -292 1236 -276
rect 1170 -346 1186 -292
rect 1220 -346 1236 -292
rect 1170 -362 1236 -346
rect 1282 -292 1356 -276
rect 1282 -346 1298 -292
rect 1340 -346 1356 -292
rect 1282 -362 1356 -346
rect 1402 -292 1468 -276
rect 1402 -346 1418 -292
rect 1452 -346 1468 -292
rect 1402 -362 1468 -346
rect 1514 -292 1588 -276
rect 1514 -346 1530 -292
rect 1572 -346 1588 -292
rect 1514 -362 1588 -346
rect 1634 -292 1700 -276
rect 1634 -346 1650 -292
rect 1684 -346 1700 -292
rect 1634 -362 1700 -346
rect 1746 -292 1820 -276
rect 1746 -346 1762 -292
rect 1804 -346 1820 -292
rect 1746 -362 1820 -346
rect 76 -426 96 -362
rect 0 -482 96 -426
<< viali >>
rect 314 268 348 302
rect 202 148 236 202
rect 546 268 580 302
rect 434 148 468 202
rect 778 268 812 302
rect 666 148 700 202
rect 1010 268 1044 302
rect 898 148 932 202
rect 1242 268 1276 302
rect 1130 148 1164 202
rect 1474 268 1508 302
rect 1362 148 1396 202
rect 1706 268 1740 302
rect 1594 148 1628 202
rect 202 -82 236 -48
rect 314 -82 348 -48
rect 434 -82 468 -48
rect 546 -82 580 -48
rect 666 -82 700 -48
rect 778 -82 812 -48
rect 898 -82 932 -48
rect 1010 -82 1044 -48
rect 1130 -82 1164 -48
rect 1242 -82 1276 -48
rect 1362 -82 1396 -48
rect 1474 -82 1508 -48
rect 1594 -82 1628 -48
rect 1706 -82 1740 -48
<< metal1 >>
rect 298 302 364 318
rect 298 268 314 302
rect 348 268 364 302
rect 186 202 252 218
rect 186 148 202 202
rect 236 148 252 202
rect 186 -48 252 148
rect 186 -82 202 -48
rect 236 -82 252 -48
rect 186 -98 252 -82
rect 298 -48 364 268
rect 530 302 596 318
rect 530 268 546 302
rect 580 268 596 302
rect 298 -82 314 -48
rect 348 -82 364 -48
rect 298 -98 364 -82
rect 418 202 484 218
rect 418 148 434 202
rect 468 148 484 202
rect 418 -48 484 148
rect 418 -82 434 -48
rect 468 -82 484 -48
rect 418 -98 484 -82
rect 530 -48 596 268
rect 762 302 828 318
rect 762 268 778 302
rect 812 268 828 302
rect 530 -82 546 -48
rect 580 -82 596 -48
rect 530 -98 596 -82
rect 650 202 716 218
rect 650 148 666 202
rect 700 148 716 202
rect 650 -48 716 148
rect 650 -82 666 -48
rect 700 -82 716 -48
rect 650 -98 716 -82
rect 762 -48 828 268
rect 994 302 1060 318
rect 994 268 1010 302
rect 1044 268 1060 302
rect 762 -82 778 -48
rect 812 -82 828 -48
rect 762 -98 828 -82
rect 882 202 948 218
rect 882 148 898 202
rect 932 148 948 202
rect 882 -48 948 148
rect 882 -82 898 -48
rect 932 -82 948 -48
rect 882 -98 948 -82
rect 994 -48 1060 268
rect 1226 302 1292 318
rect 1226 268 1242 302
rect 1276 268 1292 302
rect 994 -82 1010 -48
rect 1044 -82 1060 -48
rect 994 -98 1060 -82
rect 1114 202 1180 218
rect 1114 148 1130 202
rect 1164 148 1180 202
rect 1114 -48 1180 148
rect 1114 -82 1130 -48
rect 1164 -82 1180 -48
rect 1114 -98 1180 -82
rect 1226 -48 1292 268
rect 1458 302 1524 318
rect 1458 268 1474 302
rect 1508 268 1524 302
rect 1226 -82 1242 -48
rect 1276 -82 1292 -48
rect 1226 -98 1292 -82
rect 1346 202 1412 218
rect 1346 148 1362 202
rect 1396 148 1412 202
rect 1346 -48 1412 148
rect 1346 -82 1362 -48
rect 1396 -82 1412 -48
rect 1346 -98 1412 -82
rect 1458 -48 1524 268
rect 1690 302 1756 318
rect 1690 268 1706 302
rect 1740 268 1756 302
rect 1458 -82 1474 -48
rect 1508 -82 1524 -48
rect 1458 -98 1524 -82
rect 1578 202 1644 218
rect 1578 148 1594 202
rect 1628 148 1644 202
rect 1578 -48 1644 148
rect 1578 -82 1594 -48
rect 1628 -82 1644 -48
rect 1578 -98 1644 -82
rect 1690 -48 1756 268
rect 1690 -82 1706 -48
rect 1740 -82 1756 -48
rect 1690 -98 1756 -82
<< end >>
