magic
tech sky130A
timestamp 1739945136
<< nwell >>
rect -2 197 215 488
<< nmos >>
rect 72 65 87 115
rect 126 65 141 115
<< pmos >>
rect 72 315 87 415
rect 126 315 141 415
<< ndiff >>
rect 36 107 72 115
rect 36 73 44 107
rect 61 73 72 107
rect 36 65 72 73
rect 87 107 126 115
rect 87 73 98 107
rect 115 73 126 107
rect 87 65 126 73
rect 141 107 177 115
rect 141 73 152 107
rect 169 73 177 107
rect 141 65 177 73
<< pdiff >>
rect 36 407 72 415
rect 36 323 44 407
rect 61 323 72 407
rect 36 315 72 323
rect 87 315 126 415
rect 141 407 177 415
rect 141 323 152 407
rect 169 323 177 407
rect 141 315 177 323
<< ndiffc >>
rect 44 73 61 107
rect 98 73 115 107
rect 152 73 169 107
<< pdiffc >>
rect 44 323 61 407
rect 152 323 169 407
<< psubdiff >>
rect 0 10 12 38
rect 201 10 213 38
<< nsubdiff >>
rect 16 442 28 470
rect 185 442 197 470
<< psubdiffcont >>
rect 12 10 201 38
<< nsubdiffcont >>
rect 28 442 185 470
<< poly >>
rect 72 415 87 428
rect 126 415 141 428
rect 72 305 87 315
rect 44 290 87 305
rect 44 181 59 290
rect 126 260 141 315
rect 93 252 141 260
rect 93 235 101 252
rect 118 235 141 252
rect 93 227 141 235
rect 39 173 87 181
rect 39 156 47 173
rect 64 156 87 173
rect 39 148 87 156
rect 72 115 87 148
rect 126 115 141 227
rect 72 52 87 65
rect 126 52 141 65
<< polycont >>
rect 101 235 118 252
rect 47 156 64 173
<< locali >>
rect 0 470 213 480
rect 0 442 28 470
rect 185 442 213 470
rect 0 432 213 442
rect 36 407 69 432
rect 36 323 44 407
rect 61 323 69 407
rect 36 315 69 323
rect 144 407 177 415
rect 144 323 152 407
rect 169 323 177 407
rect 93 252 126 260
rect 93 235 101 252
rect 118 235 126 252
rect 93 227 126 235
rect 39 173 72 181
rect 144 180 177 323
rect 39 156 47 173
rect 64 156 72 173
rect 39 148 72 156
rect 90 148 177 180
rect 36 107 69 115
rect 36 73 44 107
rect 61 73 69 107
rect 36 48 69 73
rect 90 107 123 148
rect 90 73 98 107
rect 115 73 123 107
rect 90 65 123 73
rect 145 107 177 115
rect 145 73 152 107
rect 169 73 177 107
rect 145 48 177 73
rect 0 38 213 48
rect 0 10 12 38
rect 201 10 213 38
rect 0 0 213 10
<< labels >>
flabel ndiff 72 90 72 90 1 FreeSerif 8 0 0 0 S$
flabel pdiff 72 365 72 365 1 FreeSerif 8 0 0 0 S$
flabel locali 39 148 72 181 0 FreeSerif 80 0 0 0 B
port 8 nsew
flabel locali 144 148 177 315 0 FreeSerif 80 0 0 0 Y
port 5 nsew
flabel locali 0 432 213 480 0 FreeSerif 80 0 0 0 VDD!
port 2 nsew
flabel locali 0 0 213 48 0 FreeSerif 80 0 0 0 GND!
port 3 nsew
flabel ndiff 141 90 141 90 1 FreeSerif 8 0 0 0 S$
flabel pdiff 126 365 126 365 1 FreeSerif 8 0 0 0 S$
flabel locali 93 227 126 260 0 FreeSerif 80 0 0 0 A
port 4 nsew
<< end >>
