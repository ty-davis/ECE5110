magic
tech sky130A
magscale 1 2
timestamp 1745456262
<< nwell >>
rect -12 -1592 4182 -1322
rect -12 -2126 2120 -1592
<< nmos >>
rect 298 -1224 332 -1138
rect 562 -1224 596 -1138
rect 826 -1224 860 -1138
rect 1090 -1224 1124 -1138
rect 1354 -1224 1388 -1138
rect 1618 -1224 1652 -1138
rect 1882 -1224 1916 -1138
rect 2428 -1224 2462 -1138
rect 2692 -1224 2726 -1138
rect 2956 -1224 2990 -1138
rect 3220 -1224 3254 -1138
rect 3484 -1224 3518 -1138
rect 3748 -1224 3782 -1138
rect 4012 -1224 4046 -1138
rect 2352 -1808 2386 -1722
rect 2616 -1808 2650 -1722
rect 2484 -1950 2518 -1864
rect 2616 -1950 2650 -1864
rect 2880 -1808 2914 -1722
rect 2880 -1950 2914 -1864
rect 3144 -1808 3178 -1722
rect 3144 -1950 3178 -1864
rect 3408 -1808 3442 -1722
rect 3408 -1950 3442 -1864
rect 3672 -1808 3706 -1722
rect 3672 -1950 3706 -1864
rect 3936 -1808 3970 -1722
rect 3936 -1950 3970 -1864
<< pmos >>
rect 298 -1444 332 -1358
rect 562 -1444 596 -1358
rect 826 -1444 860 -1358
rect 1090 -1444 1124 -1358
rect 1354 -1444 1388 -1358
rect 1618 -1444 1652 -1358
rect 1882 -1444 1916 -1358
rect 2428 -1444 2462 -1358
rect 2692 -1444 2726 -1358
rect 2956 -1444 2990 -1358
rect 3220 -1444 3254 -1358
rect 3484 -1444 3518 -1358
rect 3748 -1444 3782 -1358
rect 4012 -1444 4046 -1358
rect 374 -1808 408 -1722
rect 374 -1950 408 -1864
rect 638 -1808 672 -1722
rect 638 -1950 672 -1864
rect 902 -1808 936 -1722
rect 902 -1950 936 -1864
rect 1166 -1808 1200 -1722
rect 1166 -1950 1200 -1864
rect 1430 -1808 1464 -1722
rect 1430 -1950 1464 -1864
rect 1694 -1808 1728 -1722
rect 1958 -1808 1992 -1722
rect 1694 -1950 1728 -1864
rect 1826 -1950 1860 -1864
<< ndiff >>
rect 226 -1154 298 -1138
rect 226 -1208 242 -1154
rect 276 -1208 298 -1154
rect 226 -1224 298 -1208
rect 332 -1154 404 -1138
rect 332 -1208 354 -1154
rect 388 -1208 404 -1154
rect 332 -1224 404 -1208
rect 490 -1154 562 -1138
rect 490 -1208 506 -1154
rect 540 -1208 562 -1154
rect 490 -1224 562 -1208
rect 596 -1154 668 -1138
rect 596 -1208 618 -1154
rect 652 -1208 668 -1154
rect 596 -1224 668 -1208
rect 754 -1154 826 -1138
rect 754 -1208 770 -1154
rect 804 -1208 826 -1154
rect 754 -1224 826 -1208
rect 860 -1154 932 -1138
rect 860 -1208 882 -1154
rect 916 -1208 932 -1154
rect 860 -1224 932 -1208
rect 1018 -1154 1090 -1138
rect 1018 -1208 1034 -1154
rect 1068 -1208 1090 -1154
rect 1018 -1224 1090 -1208
rect 1124 -1154 1196 -1138
rect 1124 -1208 1146 -1154
rect 1180 -1208 1196 -1154
rect 1124 -1224 1196 -1208
rect 1282 -1154 1354 -1138
rect 1282 -1208 1298 -1154
rect 1332 -1208 1354 -1154
rect 1282 -1224 1354 -1208
rect 1388 -1154 1460 -1138
rect 1388 -1208 1410 -1154
rect 1444 -1208 1460 -1154
rect 1388 -1224 1460 -1208
rect 1546 -1154 1618 -1138
rect 1546 -1208 1562 -1154
rect 1596 -1208 1618 -1154
rect 1546 -1224 1618 -1208
rect 1652 -1154 1724 -1138
rect 1652 -1208 1674 -1154
rect 1708 -1208 1724 -1154
rect 1652 -1224 1724 -1208
rect 1810 -1154 1882 -1138
rect 1810 -1208 1826 -1154
rect 1860 -1208 1882 -1154
rect 1810 -1224 1882 -1208
rect 1916 -1154 1988 -1138
rect 1916 -1208 1938 -1154
rect 1972 -1208 1988 -1154
rect 1916 -1224 1988 -1208
rect 2356 -1154 2428 -1138
rect 2356 -1208 2372 -1154
rect 2406 -1208 2428 -1154
rect 2356 -1224 2428 -1208
rect 2462 -1154 2534 -1138
rect 2462 -1208 2484 -1154
rect 2518 -1208 2534 -1154
rect 2462 -1224 2534 -1208
rect 2620 -1154 2692 -1138
rect 2620 -1208 2636 -1154
rect 2670 -1208 2692 -1154
rect 2620 -1224 2692 -1208
rect 2726 -1154 2798 -1138
rect 2726 -1208 2748 -1154
rect 2782 -1208 2798 -1154
rect 2726 -1224 2798 -1208
rect 2884 -1154 2956 -1138
rect 2884 -1208 2900 -1154
rect 2934 -1208 2956 -1154
rect 2884 -1224 2956 -1208
rect 2990 -1154 3062 -1138
rect 2990 -1208 3012 -1154
rect 3046 -1208 3062 -1154
rect 2990 -1224 3062 -1208
rect 3148 -1154 3220 -1138
rect 3148 -1208 3164 -1154
rect 3198 -1208 3220 -1154
rect 3148 -1224 3220 -1208
rect 3254 -1154 3326 -1138
rect 3254 -1208 3276 -1154
rect 3310 -1208 3326 -1154
rect 3254 -1224 3326 -1208
rect 3412 -1154 3484 -1138
rect 3412 -1208 3428 -1154
rect 3462 -1208 3484 -1154
rect 3412 -1224 3484 -1208
rect 3518 -1154 3590 -1138
rect 3518 -1208 3540 -1154
rect 3574 -1208 3590 -1154
rect 3518 -1224 3590 -1208
rect 3676 -1154 3748 -1138
rect 3676 -1208 3692 -1154
rect 3726 -1208 3748 -1154
rect 3676 -1224 3748 -1208
rect 3782 -1154 3854 -1138
rect 3782 -1208 3804 -1154
rect 3838 -1208 3854 -1154
rect 3782 -1224 3854 -1208
rect 3940 -1154 4012 -1138
rect 3940 -1208 3956 -1154
rect 3990 -1208 4012 -1154
rect 3940 -1224 4012 -1208
rect 4046 -1154 4118 -1138
rect 4046 -1208 4068 -1154
rect 4102 -1208 4118 -1154
rect 4046 -1224 4118 -1208
rect 2270 -1738 2352 -1722
rect 2270 -1792 2286 -1738
rect 2320 -1792 2352 -1738
rect 2270 -1808 2352 -1792
rect 2386 -1738 2468 -1722
rect 2386 -1792 2418 -1738
rect 2452 -1792 2468 -1738
rect 2386 -1808 2468 -1792
rect 2534 -1738 2616 -1722
rect 2534 -1792 2550 -1738
rect 2584 -1792 2616 -1738
rect 2534 -1808 2616 -1792
rect 2650 -1738 2732 -1722
rect 2650 -1792 2682 -1738
rect 2716 -1792 2732 -1738
rect 2650 -1808 2732 -1792
rect 2402 -1880 2484 -1864
rect 2402 -1934 2418 -1880
rect 2452 -1934 2484 -1880
rect 2402 -1950 2484 -1934
rect 2518 -1880 2616 -1864
rect 2518 -1934 2550 -1880
rect 2584 -1934 2616 -1880
rect 2518 -1950 2616 -1934
rect 2650 -1880 2732 -1864
rect 2650 -1934 2682 -1880
rect 2716 -1934 2732 -1880
rect 2650 -1950 2732 -1934
rect 2798 -1738 2880 -1722
rect 2798 -1792 2814 -1738
rect 2848 -1792 2880 -1738
rect 2798 -1808 2880 -1792
rect 2914 -1738 2996 -1722
rect 2914 -1792 2946 -1738
rect 2980 -1792 2996 -1738
rect 2914 -1808 2996 -1792
rect 2798 -1880 2880 -1864
rect 2798 -1934 2814 -1880
rect 2848 -1934 2880 -1880
rect 2798 -1950 2880 -1934
rect 2914 -1880 2996 -1864
rect 2914 -1934 2946 -1880
rect 2980 -1934 2996 -1880
rect 2914 -1950 2996 -1934
rect 3062 -1738 3144 -1722
rect 3062 -1792 3078 -1738
rect 3112 -1792 3144 -1738
rect 3062 -1808 3144 -1792
rect 3178 -1738 3260 -1722
rect 3178 -1792 3210 -1738
rect 3244 -1792 3260 -1738
rect 3178 -1808 3260 -1792
rect 3062 -1880 3144 -1864
rect 3062 -1934 3078 -1880
rect 3112 -1934 3144 -1880
rect 3062 -1950 3144 -1934
rect 3178 -1880 3260 -1864
rect 3178 -1934 3210 -1880
rect 3244 -1934 3260 -1880
rect 3178 -1950 3260 -1934
rect 3326 -1738 3408 -1722
rect 3326 -1792 3342 -1738
rect 3376 -1792 3408 -1738
rect 3326 -1808 3408 -1792
rect 3442 -1738 3524 -1722
rect 3442 -1792 3474 -1738
rect 3508 -1792 3524 -1738
rect 3442 -1808 3524 -1792
rect 3326 -1880 3408 -1864
rect 3326 -1934 3342 -1880
rect 3376 -1934 3408 -1880
rect 3326 -1950 3408 -1934
rect 3442 -1880 3524 -1864
rect 3442 -1934 3474 -1880
rect 3508 -1934 3524 -1880
rect 3442 -1950 3524 -1934
rect 3590 -1738 3672 -1722
rect 3590 -1792 3606 -1738
rect 3640 -1792 3672 -1738
rect 3590 -1808 3672 -1792
rect 3706 -1738 3788 -1722
rect 3706 -1792 3738 -1738
rect 3772 -1792 3788 -1738
rect 3706 -1808 3788 -1792
rect 3590 -1880 3672 -1864
rect 3590 -1934 3606 -1880
rect 3640 -1934 3672 -1880
rect 3590 -1950 3672 -1934
rect 3706 -1880 3788 -1864
rect 3706 -1934 3738 -1880
rect 3772 -1934 3788 -1880
rect 3706 -1950 3788 -1934
rect 3854 -1738 3936 -1722
rect 3854 -1792 3870 -1738
rect 3904 -1792 3936 -1738
rect 3854 -1808 3936 -1792
rect 3970 -1738 4052 -1722
rect 3970 -1792 4002 -1738
rect 4036 -1792 4052 -1738
rect 3970 -1808 4052 -1792
rect 3854 -1880 3936 -1864
rect 3854 -1934 3870 -1880
rect 3904 -1934 3936 -1880
rect 3854 -1950 3936 -1934
rect 3970 -1880 4052 -1864
rect 3970 -1934 4002 -1880
rect 4036 -1934 4052 -1880
rect 3970 -1950 4052 -1934
<< pdiff >>
rect 226 -1374 298 -1358
rect 226 -1428 242 -1374
rect 276 -1428 298 -1374
rect 226 -1444 298 -1428
rect 332 -1374 404 -1358
rect 332 -1428 354 -1374
rect 388 -1428 404 -1374
rect 332 -1444 404 -1428
rect 490 -1374 562 -1358
rect 490 -1428 506 -1374
rect 540 -1428 562 -1374
rect 490 -1444 562 -1428
rect 596 -1374 668 -1358
rect 596 -1428 618 -1374
rect 652 -1428 668 -1374
rect 596 -1444 668 -1428
rect 754 -1374 826 -1358
rect 754 -1428 770 -1374
rect 804 -1428 826 -1374
rect 754 -1444 826 -1428
rect 860 -1374 932 -1358
rect 860 -1428 882 -1374
rect 916 -1428 932 -1374
rect 860 -1444 932 -1428
rect 1018 -1374 1090 -1358
rect 1018 -1428 1034 -1374
rect 1068 -1428 1090 -1374
rect 1018 -1444 1090 -1428
rect 1124 -1374 1196 -1358
rect 1124 -1428 1146 -1374
rect 1180 -1428 1196 -1374
rect 1124 -1444 1196 -1428
rect 1282 -1374 1354 -1358
rect 1282 -1428 1298 -1374
rect 1332 -1428 1354 -1374
rect 1282 -1444 1354 -1428
rect 1388 -1374 1460 -1358
rect 1388 -1428 1410 -1374
rect 1444 -1428 1460 -1374
rect 1388 -1444 1460 -1428
rect 1546 -1374 1618 -1358
rect 1546 -1428 1562 -1374
rect 1596 -1428 1618 -1374
rect 1546 -1444 1618 -1428
rect 1652 -1374 1724 -1358
rect 1652 -1428 1674 -1374
rect 1708 -1428 1724 -1374
rect 1652 -1444 1724 -1428
rect 1810 -1374 1882 -1358
rect 1810 -1428 1826 -1374
rect 1860 -1428 1882 -1374
rect 1810 -1444 1882 -1428
rect 1916 -1374 1988 -1358
rect 1916 -1428 1938 -1374
rect 1972 -1428 1988 -1374
rect 1916 -1444 1988 -1428
rect 2356 -1374 2428 -1358
rect 2356 -1428 2372 -1374
rect 2406 -1428 2428 -1374
rect 2356 -1444 2428 -1428
rect 2462 -1374 2534 -1358
rect 2462 -1428 2484 -1374
rect 2518 -1428 2534 -1374
rect 2462 -1444 2534 -1428
rect 2620 -1374 2692 -1358
rect 2620 -1428 2636 -1374
rect 2670 -1428 2692 -1374
rect 2620 -1444 2692 -1428
rect 2726 -1374 2798 -1358
rect 2726 -1428 2748 -1374
rect 2782 -1428 2798 -1374
rect 2726 -1444 2798 -1428
rect 2884 -1374 2956 -1358
rect 2884 -1428 2900 -1374
rect 2934 -1428 2956 -1374
rect 2884 -1444 2956 -1428
rect 2990 -1374 3062 -1358
rect 2990 -1428 3012 -1374
rect 3046 -1428 3062 -1374
rect 2990 -1444 3062 -1428
rect 3148 -1374 3220 -1358
rect 3148 -1428 3164 -1374
rect 3198 -1428 3220 -1374
rect 3148 -1444 3220 -1428
rect 3254 -1374 3326 -1358
rect 3254 -1428 3276 -1374
rect 3310 -1428 3326 -1374
rect 3254 -1444 3326 -1428
rect 3412 -1374 3484 -1358
rect 3412 -1428 3428 -1374
rect 3462 -1428 3484 -1374
rect 3412 -1444 3484 -1428
rect 3518 -1374 3590 -1358
rect 3518 -1428 3540 -1374
rect 3574 -1428 3590 -1374
rect 3518 -1444 3590 -1428
rect 3676 -1374 3748 -1358
rect 3676 -1428 3692 -1374
rect 3726 -1428 3748 -1374
rect 3676 -1444 3748 -1428
rect 3782 -1374 3854 -1358
rect 3782 -1428 3804 -1374
rect 3838 -1428 3854 -1374
rect 3782 -1444 3854 -1428
rect 3940 -1374 4012 -1358
rect 3940 -1428 3956 -1374
rect 3990 -1428 4012 -1374
rect 3940 -1444 4012 -1428
rect 4046 -1374 4118 -1358
rect 4046 -1428 4068 -1374
rect 4102 -1428 4118 -1374
rect 4046 -1444 4118 -1428
rect 160 -1738 226 -1722
rect 160 -1792 176 -1738
rect 210 -1792 226 -1738
rect 160 -1808 226 -1792
rect 160 -1880 226 -1864
rect 160 -1934 176 -1880
rect 210 -1934 226 -1880
rect 160 -1950 226 -1934
rect 292 -1738 374 -1722
rect 292 -1792 308 -1738
rect 342 -1792 374 -1738
rect 292 -1808 374 -1792
rect 408 -1738 490 -1722
rect 408 -1792 440 -1738
rect 474 -1792 490 -1738
rect 408 -1808 490 -1792
rect 292 -1880 374 -1864
rect 292 -1934 308 -1880
rect 342 -1934 374 -1880
rect 292 -1950 374 -1934
rect 408 -1880 490 -1864
rect 408 -1934 440 -1880
rect 474 -1934 490 -1880
rect 408 -1950 490 -1934
rect 556 -1738 638 -1722
rect 556 -1792 572 -1738
rect 606 -1792 638 -1738
rect 556 -1808 638 -1792
rect 672 -1738 754 -1722
rect 672 -1792 704 -1738
rect 738 -1792 754 -1738
rect 672 -1808 754 -1792
rect 556 -1880 638 -1864
rect 556 -1934 572 -1880
rect 606 -1934 638 -1880
rect 556 -1950 638 -1934
rect 672 -1880 754 -1864
rect 672 -1934 704 -1880
rect 738 -1934 754 -1880
rect 672 -1950 754 -1934
rect 820 -1738 902 -1722
rect 820 -1792 836 -1738
rect 870 -1792 902 -1738
rect 820 -1808 902 -1792
rect 936 -1738 1018 -1722
rect 936 -1792 968 -1738
rect 1002 -1792 1018 -1738
rect 936 -1808 1018 -1792
rect 820 -1880 902 -1864
rect 820 -1934 836 -1880
rect 870 -1934 902 -1880
rect 820 -1950 902 -1934
rect 936 -1880 1018 -1864
rect 936 -1934 968 -1880
rect 1002 -1934 1018 -1880
rect 936 -1950 1018 -1934
rect 1084 -1738 1166 -1722
rect 1084 -1792 1100 -1738
rect 1134 -1792 1166 -1738
rect 1084 -1808 1166 -1792
rect 1200 -1738 1282 -1722
rect 1200 -1792 1232 -1738
rect 1266 -1792 1282 -1738
rect 1200 -1808 1282 -1792
rect 1084 -1880 1166 -1864
rect 1084 -1934 1100 -1880
rect 1134 -1934 1166 -1880
rect 1084 -1950 1166 -1934
rect 1200 -1880 1282 -1864
rect 1200 -1934 1232 -1880
rect 1266 -1934 1282 -1880
rect 1200 -1950 1282 -1934
rect 1348 -1738 1430 -1722
rect 1348 -1792 1364 -1738
rect 1398 -1792 1430 -1738
rect 1348 -1808 1430 -1792
rect 1464 -1738 1546 -1722
rect 1464 -1792 1496 -1738
rect 1530 -1792 1546 -1738
rect 1464 -1808 1546 -1792
rect 1348 -1880 1430 -1864
rect 1348 -1934 1364 -1880
rect 1398 -1934 1430 -1880
rect 1348 -1950 1430 -1934
rect 1464 -1880 1546 -1864
rect 1464 -1934 1496 -1880
rect 1530 -1934 1546 -1880
rect 1464 -1950 1546 -1934
rect 1612 -1738 1694 -1722
rect 1612 -1792 1628 -1738
rect 1662 -1792 1694 -1738
rect 1612 -1808 1694 -1792
rect 1728 -1738 1810 -1722
rect 1728 -1792 1760 -1738
rect 1794 -1792 1810 -1738
rect 1728 -1808 1810 -1792
rect 1876 -1738 1958 -1722
rect 1876 -1792 1892 -1738
rect 1926 -1792 1958 -1738
rect 1876 -1808 1958 -1792
rect 1992 -1738 2074 -1722
rect 1992 -1792 2024 -1738
rect 2058 -1792 2074 -1738
rect 1992 -1808 2074 -1792
rect 1612 -1880 1694 -1864
rect 1612 -1934 1628 -1880
rect 1662 -1934 1694 -1880
rect 1612 -1950 1694 -1934
rect 1728 -1880 1826 -1864
rect 1728 -1934 1760 -1880
rect 1794 -1934 1826 -1880
rect 1728 -1950 1826 -1934
rect 1860 -1880 1942 -1864
rect 1860 -1934 1892 -1880
rect 1926 -1934 1942 -1880
rect 1860 -1950 1942 -1934
rect 2008 -1880 2074 -1864
rect 2008 -1934 2024 -1880
rect 2058 -1934 2074 -1880
rect 2008 -1950 2074 -1934
<< ndiffc >>
rect 242 -1208 276 -1154
rect 354 -1208 388 -1154
rect 506 -1208 540 -1154
rect 618 -1208 652 -1154
rect 770 -1208 804 -1154
rect 882 -1208 916 -1154
rect 1034 -1208 1068 -1154
rect 1146 -1208 1180 -1154
rect 1298 -1208 1332 -1154
rect 1410 -1208 1444 -1154
rect 1562 -1208 1596 -1154
rect 1674 -1208 1708 -1154
rect 1826 -1208 1860 -1154
rect 1938 -1208 1972 -1154
rect 2372 -1208 2406 -1154
rect 2484 -1208 2518 -1154
rect 2636 -1208 2670 -1154
rect 2748 -1208 2782 -1154
rect 2900 -1208 2934 -1154
rect 3012 -1208 3046 -1154
rect 3164 -1208 3198 -1154
rect 3276 -1208 3310 -1154
rect 3428 -1208 3462 -1154
rect 3540 -1208 3574 -1154
rect 3692 -1208 3726 -1154
rect 3804 -1208 3838 -1154
rect 3956 -1208 3990 -1154
rect 4068 -1208 4102 -1154
rect 2286 -1792 2320 -1738
rect 2418 -1792 2452 -1738
rect 2550 -1792 2584 -1738
rect 2682 -1792 2716 -1738
rect 2418 -1934 2452 -1880
rect 2550 -1934 2584 -1880
rect 2682 -1934 2716 -1880
rect 2814 -1792 2848 -1738
rect 2946 -1792 2980 -1738
rect 2814 -1934 2848 -1880
rect 2946 -1934 2980 -1880
rect 3078 -1792 3112 -1738
rect 3210 -1792 3244 -1738
rect 3078 -1934 3112 -1880
rect 3210 -1934 3244 -1880
rect 3342 -1792 3376 -1738
rect 3474 -1792 3508 -1738
rect 3342 -1934 3376 -1880
rect 3474 -1934 3508 -1880
rect 3606 -1792 3640 -1738
rect 3738 -1792 3772 -1738
rect 3606 -1934 3640 -1880
rect 3738 -1934 3772 -1880
rect 3870 -1792 3904 -1738
rect 4002 -1792 4036 -1738
rect 3870 -1934 3904 -1880
rect 4002 -1934 4036 -1880
<< pdiffc >>
rect 242 -1428 276 -1374
rect 354 -1428 388 -1374
rect 506 -1428 540 -1374
rect 618 -1428 652 -1374
rect 770 -1428 804 -1374
rect 882 -1428 916 -1374
rect 1034 -1428 1068 -1374
rect 1146 -1428 1180 -1374
rect 1298 -1428 1332 -1374
rect 1410 -1428 1444 -1374
rect 1562 -1428 1596 -1374
rect 1674 -1428 1708 -1374
rect 1826 -1428 1860 -1374
rect 1938 -1428 1972 -1374
rect 2372 -1428 2406 -1374
rect 2484 -1428 2518 -1374
rect 2636 -1428 2670 -1374
rect 2748 -1428 2782 -1374
rect 2900 -1428 2934 -1374
rect 3012 -1428 3046 -1374
rect 3164 -1428 3198 -1374
rect 3276 -1428 3310 -1374
rect 3428 -1428 3462 -1374
rect 3540 -1428 3574 -1374
rect 3692 -1428 3726 -1374
rect 3804 -1428 3838 -1374
rect 3956 -1428 3990 -1374
rect 4068 -1428 4102 -1374
rect 176 -1792 210 -1738
rect 176 -1934 210 -1880
rect 308 -1792 342 -1738
rect 440 -1792 474 -1738
rect 308 -1934 342 -1880
rect 440 -1934 474 -1880
rect 572 -1792 606 -1738
rect 704 -1792 738 -1738
rect 572 -1934 606 -1880
rect 704 -1934 738 -1880
rect 836 -1792 870 -1738
rect 968 -1792 1002 -1738
rect 836 -1934 870 -1880
rect 968 -1934 1002 -1880
rect 1100 -1792 1134 -1738
rect 1232 -1792 1266 -1738
rect 1100 -1934 1134 -1880
rect 1232 -1934 1266 -1880
rect 1364 -1792 1398 -1738
rect 1496 -1792 1530 -1738
rect 1364 -1934 1398 -1880
rect 1496 -1934 1530 -1880
rect 1628 -1792 1662 -1738
rect 1760 -1792 1794 -1738
rect 1892 -1792 1926 -1738
rect 2024 -1792 2058 -1738
rect 1628 -1934 1662 -1880
rect 1760 -1934 1794 -1880
rect 1892 -1934 1926 -1880
rect 2024 -1934 2058 -1880
<< psubdiff >>
rect 48 -1084 72 -1028
rect 4090 -1084 4114 -1028
rect 2162 -2200 2186 -2144
rect 4090 -2200 4114 -2144
<< nsubdiff >>
rect 48 -1554 72 -1498
rect 4122 -1554 4146 -1498
rect 44 -1632 100 -1608
rect 44 -2060 46 -1632
rect 44 -2084 100 -2060
<< psubdiffcont >>
rect 72 -1084 4090 -1028
rect 2186 -2200 4090 -2144
<< nsubdiffcont >>
rect 72 -1554 4122 -1498
rect 46 -2060 100 -1632
<< poly >>
rect 298 -1138 332 -1112
rect 562 -1138 596 -1112
rect 826 -1138 860 -1112
rect 1090 -1138 1124 -1112
rect 1354 -1138 1388 -1112
rect 1618 -1138 1652 -1112
rect 1882 -1138 1916 -1112
rect 2428 -1138 2462 -1112
rect 2692 -1138 2726 -1112
rect 2956 -1138 2990 -1112
rect 3220 -1138 3254 -1112
rect 3484 -1138 3518 -1112
rect 3748 -1138 3782 -1112
rect 4012 -1138 4046 -1112
rect 298 -1258 332 -1224
rect 562 -1258 596 -1224
rect 826 -1258 860 -1224
rect 1090 -1258 1124 -1224
rect 1354 -1258 1388 -1224
rect 1618 -1258 1652 -1224
rect 1882 -1258 1916 -1224
rect 2428 -1258 2462 -1224
rect 2692 -1258 2726 -1224
rect 2956 -1258 2990 -1224
rect 3220 -1258 3254 -1224
rect 3484 -1258 3518 -1224
rect 3748 -1258 3782 -1224
rect 4012 -1258 4046 -1224
rect 298 -1274 404 -1258
rect 298 -1308 354 -1274
rect 388 -1308 404 -1274
rect 298 -1324 404 -1308
rect 562 -1274 668 -1258
rect 562 -1308 618 -1274
rect 652 -1308 668 -1274
rect 562 -1324 668 -1308
rect 826 -1274 932 -1258
rect 826 -1308 882 -1274
rect 916 -1308 932 -1274
rect 826 -1324 932 -1308
rect 1090 -1274 1196 -1258
rect 1090 -1308 1146 -1274
rect 1180 -1308 1196 -1274
rect 1090 -1324 1196 -1308
rect 1354 -1274 1460 -1258
rect 1354 -1308 1410 -1274
rect 1444 -1308 1460 -1274
rect 1354 -1324 1460 -1308
rect 1618 -1274 1724 -1258
rect 1618 -1308 1674 -1274
rect 1708 -1308 1724 -1274
rect 1618 -1324 1724 -1308
rect 1882 -1274 1988 -1258
rect 1882 -1308 1938 -1274
rect 1972 -1308 1988 -1274
rect 1882 -1324 1988 -1308
rect 2356 -1274 2462 -1258
rect 2356 -1308 2372 -1274
rect 2406 -1308 2462 -1274
rect 2356 -1324 2462 -1308
rect 2620 -1274 2726 -1258
rect 2620 -1308 2636 -1274
rect 2670 -1308 2726 -1274
rect 2620 -1324 2726 -1308
rect 2884 -1274 2990 -1258
rect 2884 -1308 2900 -1274
rect 2934 -1308 2990 -1274
rect 2884 -1324 2990 -1308
rect 3148 -1274 3254 -1258
rect 3148 -1308 3164 -1274
rect 3198 -1308 3254 -1274
rect 3148 -1324 3254 -1308
rect 3412 -1274 3518 -1258
rect 3412 -1308 3428 -1274
rect 3462 -1308 3518 -1274
rect 3412 -1324 3518 -1308
rect 3676 -1274 3782 -1258
rect 3676 -1308 3692 -1274
rect 3726 -1308 3782 -1274
rect 3676 -1324 3782 -1308
rect 3940 -1274 4046 -1258
rect 3940 -1308 3956 -1274
rect 3990 -1308 4046 -1274
rect 3940 -1324 4046 -1308
rect 298 -1358 332 -1324
rect 562 -1358 596 -1324
rect 826 -1358 860 -1324
rect 1090 -1358 1124 -1324
rect 1354 -1358 1388 -1324
rect 1618 -1358 1652 -1324
rect 1882 -1358 1916 -1324
rect 2428 -1358 2462 -1324
rect 2692 -1358 2726 -1324
rect 2956 -1358 2990 -1324
rect 3220 -1358 3254 -1324
rect 3484 -1358 3518 -1324
rect 3748 -1358 3782 -1324
rect 4012 -1358 4046 -1324
rect 298 -1470 332 -1444
rect 562 -1470 596 -1444
rect 826 -1470 860 -1444
rect 1090 -1470 1124 -1444
rect 1354 -1470 1388 -1444
rect 1618 -1470 1652 -1444
rect 1882 -1470 1916 -1444
rect 2428 -1470 2462 -1444
rect 2692 -1470 2726 -1444
rect 2956 -1470 2990 -1444
rect 3220 -1470 3254 -1444
rect 3484 -1470 3518 -1444
rect 3748 -1470 3782 -1444
rect 4012 -1470 4046 -1444
rect 226 -1624 292 -1608
rect 226 -1658 242 -1624
rect 276 -1658 292 -1624
rect 226 -1674 292 -1658
rect 358 -1624 424 -1608
rect 358 -1658 374 -1624
rect 408 -1658 424 -1624
rect 358 -1674 424 -1658
rect 490 -1624 556 -1608
rect 490 -1658 506 -1624
rect 540 -1658 556 -1624
rect 490 -1674 556 -1658
rect 622 -1624 688 -1608
rect 622 -1658 638 -1624
rect 672 -1658 688 -1624
rect 622 -1674 688 -1658
rect 754 -1624 820 -1608
rect 754 -1658 770 -1624
rect 804 -1658 820 -1624
rect 754 -1674 820 -1658
rect 886 -1624 952 -1608
rect 886 -1658 902 -1624
rect 936 -1658 952 -1624
rect 886 -1674 952 -1658
rect 1018 -1624 1084 -1608
rect 1018 -1658 1034 -1624
rect 1068 -1658 1084 -1624
rect 1018 -1674 1084 -1658
rect 1150 -1624 1216 -1608
rect 1150 -1658 1166 -1624
rect 1200 -1658 1216 -1624
rect 1150 -1674 1216 -1658
rect 1282 -1624 1348 -1608
rect 1282 -1658 1298 -1624
rect 1332 -1658 1348 -1624
rect 1282 -1674 1348 -1658
rect 1414 -1624 1480 -1608
rect 1414 -1658 1430 -1624
rect 1464 -1658 1480 -1624
rect 1414 -1674 1480 -1658
rect 1546 -1624 1612 -1608
rect 1546 -1658 1562 -1624
rect 1596 -1658 1612 -1624
rect 1546 -1674 1612 -1658
rect 1678 -1624 1744 -1608
rect 1678 -1658 1694 -1624
rect 1728 -1658 1744 -1624
rect 1678 -1674 1744 -1658
rect 1810 -1624 1876 -1608
rect 1810 -1658 1826 -1624
rect 1860 -1658 1876 -1624
rect 1810 -1674 1876 -1658
rect 1942 -1624 2008 -1608
rect 1942 -1658 1958 -1624
rect 1992 -1658 2008 -1624
rect 1942 -1674 2008 -1658
rect 2336 -1624 2402 -1608
rect 2336 -1658 2352 -1624
rect 2386 -1658 2402 -1624
rect 2336 -1674 2402 -1658
rect 2468 -1624 2534 -1608
rect 2468 -1658 2484 -1624
rect 2518 -1658 2534 -1624
rect 2468 -1674 2534 -1658
rect 2600 -1624 2666 -1608
rect 2600 -1658 2616 -1624
rect 2650 -1658 2666 -1624
rect 2600 -1674 2666 -1658
rect 2732 -1624 2798 -1608
rect 2732 -1658 2748 -1624
rect 2782 -1658 2798 -1624
rect 2732 -1674 2798 -1658
rect 2864 -1624 2930 -1608
rect 2864 -1658 2880 -1624
rect 2914 -1658 2930 -1624
rect 2864 -1674 2930 -1658
rect 2996 -1624 3062 -1608
rect 2996 -1658 3012 -1624
rect 3046 -1658 3062 -1624
rect 2996 -1674 3062 -1658
rect 3128 -1624 3194 -1608
rect 3128 -1658 3144 -1624
rect 3178 -1658 3194 -1624
rect 3128 -1674 3194 -1658
rect 3260 -1624 3326 -1608
rect 3260 -1658 3276 -1624
rect 3310 -1658 3326 -1624
rect 3260 -1674 3326 -1658
rect 3392 -1624 3458 -1608
rect 3392 -1658 3408 -1624
rect 3442 -1658 3458 -1624
rect 3392 -1674 3458 -1658
rect 3524 -1624 3590 -1608
rect 3524 -1658 3540 -1624
rect 3574 -1658 3590 -1624
rect 3524 -1674 3590 -1658
rect 3656 -1624 3722 -1608
rect 3656 -1658 3672 -1624
rect 3706 -1658 3722 -1624
rect 3656 -1674 3722 -1658
rect 3788 -1624 3854 -1608
rect 3788 -1658 3804 -1624
rect 3838 -1658 3854 -1624
rect 3788 -1674 3854 -1658
rect 3920 -1624 3986 -1608
rect 3920 -1658 3936 -1624
rect 3970 -1658 3986 -1624
rect 3920 -1674 3986 -1658
rect 4052 -1624 4118 -1608
rect 4052 -1658 4068 -1624
rect 4102 -1658 4118 -1624
rect 4052 -1674 4118 -1658
rect 242 -1976 276 -1674
rect 374 -1722 408 -1674
rect 374 -1864 408 -1808
rect 374 -1976 408 -1950
rect 506 -1976 540 -1674
rect 638 -1722 672 -1674
rect 638 -1864 672 -1808
rect 638 -1976 672 -1950
rect 770 -1976 804 -1674
rect 902 -1722 936 -1674
rect 902 -1864 936 -1808
rect 902 -1976 936 -1950
rect 1034 -1976 1068 -1674
rect 1166 -1722 1200 -1674
rect 1166 -1864 1200 -1808
rect 1166 -1976 1200 -1950
rect 1298 -1976 1332 -1674
rect 1430 -1722 1464 -1674
rect 1430 -1864 1464 -1808
rect 1430 -1976 1464 -1950
rect 1562 -1976 1596 -1674
rect 1694 -1722 1728 -1674
rect 1694 -1864 1728 -1808
rect 1826 -1864 1860 -1674
rect 1958 -1722 1992 -1674
rect 2352 -1722 2386 -1674
rect 1694 -1976 1728 -1950
rect 1826 -1976 1860 -1950
rect 1958 -1976 1992 -1808
rect 2352 -1976 2386 -1808
rect 2484 -1864 2518 -1674
rect 2616 -1722 2650 -1674
rect 2616 -1864 2650 -1808
rect 2484 -1976 2518 -1950
rect 2616 -1976 2650 -1950
rect 2748 -1976 2782 -1674
rect 2880 -1722 2914 -1674
rect 2880 -1864 2914 -1808
rect 2880 -1976 2914 -1950
rect 3012 -1976 3046 -1674
rect 3144 -1722 3178 -1674
rect 3144 -1864 3178 -1808
rect 3144 -1976 3178 -1950
rect 3276 -1976 3310 -1674
rect 3408 -1722 3442 -1674
rect 3408 -1864 3442 -1808
rect 3408 -1976 3442 -1950
rect 3540 -1976 3574 -1674
rect 3672 -1722 3706 -1674
rect 3672 -1864 3706 -1808
rect 3672 -1976 3706 -1950
rect 3804 -1976 3838 -1674
rect 3936 -1722 3970 -1674
rect 3936 -1864 3970 -1808
rect 3936 -1976 3970 -1950
rect 4068 -1976 4102 -1674
<< polycont >>
rect 354 -1308 388 -1274
rect 618 -1308 652 -1274
rect 882 -1308 916 -1274
rect 1146 -1308 1180 -1274
rect 1410 -1308 1444 -1274
rect 1674 -1308 1708 -1274
rect 1938 -1308 1972 -1274
rect 2372 -1308 2406 -1274
rect 2636 -1308 2670 -1274
rect 2900 -1308 2934 -1274
rect 3164 -1308 3198 -1274
rect 3428 -1308 3462 -1274
rect 3692 -1308 3726 -1274
rect 3956 -1308 3990 -1274
rect 242 -1658 276 -1624
rect 374 -1658 408 -1624
rect 506 -1658 540 -1624
rect 638 -1658 672 -1624
rect 770 -1658 804 -1624
rect 902 -1658 936 -1624
rect 1034 -1658 1068 -1624
rect 1166 -1658 1200 -1624
rect 1298 -1658 1332 -1624
rect 1430 -1658 1464 -1624
rect 1562 -1658 1596 -1624
rect 1694 -1658 1728 -1624
rect 1826 -1658 1860 -1624
rect 1958 -1658 1992 -1624
rect 2352 -1658 2386 -1624
rect 2484 -1658 2518 -1624
rect 2616 -1658 2650 -1624
rect 2748 -1658 2782 -1624
rect 2880 -1658 2914 -1624
rect 3012 -1658 3046 -1624
rect 3144 -1658 3178 -1624
rect 3276 -1658 3310 -1624
rect 3408 -1658 3442 -1624
rect 3540 -1658 3574 -1624
rect 3672 -1658 3706 -1624
rect 3804 -1658 3838 -1624
rect 3936 -1658 3970 -1624
rect 4068 -1658 4102 -1624
<< locali >>
rect 24 -1028 4294 -1008
rect 24 -1084 72 -1028
rect 4090 -1084 4294 -1028
rect 24 -1104 4294 -1084
rect 226 -1154 292 -1138
rect 226 -1208 242 -1154
rect 276 -1208 292 -1154
rect 226 -1374 292 -1208
rect 338 -1154 404 -1104
rect 338 -1208 354 -1154
rect 388 -1208 404 -1154
rect 338 -1224 404 -1208
rect 490 -1154 556 -1138
rect 490 -1208 506 -1154
rect 540 -1208 556 -1154
rect 332 -1274 404 -1258
rect 332 -1308 354 -1274
rect 388 -1308 404 -1274
rect 332 -1324 404 -1308
rect 226 -1428 242 -1374
rect 276 -1428 292 -1374
rect 226 -1444 292 -1428
rect 338 -1374 404 -1358
rect 338 -1428 354 -1374
rect 388 -1428 404 -1374
rect 338 -1478 404 -1428
rect 490 -1374 556 -1208
rect 602 -1154 668 -1104
rect 602 -1208 618 -1154
rect 652 -1208 668 -1154
rect 602 -1224 668 -1208
rect 754 -1154 820 -1138
rect 754 -1208 770 -1154
rect 804 -1208 820 -1154
rect 596 -1274 668 -1258
rect 596 -1308 618 -1274
rect 652 -1308 668 -1274
rect 596 -1324 668 -1308
rect 490 -1428 506 -1374
rect 540 -1428 556 -1374
rect 490 -1444 556 -1428
rect 602 -1374 668 -1358
rect 602 -1428 618 -1374
rect 652 -1428 668 -1374
rect 602 -1478 668 -1428
rect 754 -1374 820 -1208
rect 866 -1154 932 -1104
rect 866 -1208 882 -1154
rect 916 -1208 932 -1154
rect 866 -1224 932 -1208
rect 1018 -1154 1084 -1138
rect 1018 -1208 1034 -1154
rect 1068 -1208 1084 -1154
rect 860 -1274 932 -1258
rect 860 -1308 882 -1274
rect 916 -1308 932 -1274
rect 860 -1324 932 -1308
rect 754 -1428 770 -1374
rect 804 -1428 820 -1374
rect 754 -1444 820 -1428
rect 866 -1374 932 -1358
rect 866 -1428 882 -1374
rect 916 -1428 932 -1374
rect 866 -1478 932 -1428
rect 1018 -1374 1084 -1208
rect 1130 -1154 1196 -1104
rect 1130 -1208 1146 -1154
rect 1180 -1208 1196 -1154
rect 1130 -1224 1196 -1208
rect 1282 -1154 1348 -1138
rect 1282 -1208 1298 -1154
rect 1332 -1208 1348 -1154
rect 1124 -1274 1196 -1258
rect 1124 -1308 1146 -1274
rect 1180 -1308 1196 -1274
rect 1124 -1324 1196 -1308
rect 1018 -1428 1034 -1374
rect 1068 -1428 1084 -1374
rect 1018 -1444 1084 -1428
rect 1130 -1374 1196 -1358
rect 1130 -1428 1146 -1374
rect 1180 -1428 1196 -1374
rect 1130 -1478 1196 -1428
rect 1282 -1374 1348 -1208
rect 1394 -1154 1460 -1104
rect 1394 -1208 1410 -1154
rect 1444 -1208 1460 -1154
rect 1394 -1224 1460 -1208
rect 1546 -1154 1612 -1138
rect 1546 -1208 1562 -1154
rect 1596 -1208 1612 -1154
rect 1388 -1274 1460 -1258
rect 1388 -1308 1410 -1274
rect 1444 -1308 1460 -1274
rect 1388 -1324 1460 -1308
rect 1282 -1428 1298 -1374
rect 1332 -1428 1348 -1374
rect 1282 -1444 1348 -1428
rect 1394 -1374 1460 -1358
rect 1394 -1428 1410 -1374
rect 1444 -1428 1460 -1374
rect 1394 -1478 1460 -1428
rect 1546 -1374 1612 -1208
rect 1658 -1154 1724 -1104
rect 1658 -1208 1674 -1154
rect 1708 -1208 1724 -1154
rect 1658 -1224 1724 -1208
rect 1810 -1154 1876 -1138
rect 1810 -1208 1826 -1154
rect 1860 -1208 1876 -1154
rect 1652 -1274 1724 -1258
rect 1652 -1308 1674 -1274
rect 1708 -1308 1724 -1274
rect 1652 -1324 1724 -1308
rect 1546 -1428 1562 -1374
rect 1596 -1428 1612 -1374
rect 1546 -1444 1612 -1428
rect 1658 -1374 1724 -1358
rect 1658 -1428 1674 -1374
rect 1708 -1428 1724 -1374
rect 1658 -1478 1724 -1428
rect 1810 -1374 1876 -1208
rect 1922 -1154 1988 -1104
rect 1922 -1208 1938 -1154
rect 1972 -1208 1988 -1154
rect 1922 -1224 1988 -1208
rect 2356 -1154 2422 -1104
rect 2356 -1208 2372 -1154
rect 2406 -1208 2422 -1154
rect 2356 -1224 2422 -1208
rect 2468 -1154 2534 -1138
rect 2468 -1208 2484 -1154
rect 2518 -1208 2534 -1154
rect 1916 -1274 1988 -1258
rect 1916 -1308 1938 -1274
rect 1972 -1308 1988 -1274
rect 1916 -1324 1988 -1308
rect 2356 -1274 2428 -1258
rect 2356 -1308 2372 -1274
rect 2406 -1308 2428 -1274
rect 2356 -1324 2428 -1308
rect 1810 -1428 1826 -1374
rect 1860 -1428 1876 -1374
rect 1810 -1444 1876 -1428
rect 1922 -1374 1988 -1358
rect 1922 -1428 1938 -1374
rect 1972 -1428 1988 -1374
rect 1922 -1478 1988 -1428
rect 2356 -1374 2422 -1358
rect 2356 -1428 2372 -1374
rect 2406 -1428 2422 -1374
rect 2356 -1478 2422 -1428
rect 2468 -1374 2534 -1208
rect 2620 -1154 2686 -1104
rect 2620 -1208 2636 -1154
rect 2670 -1208 2686 -1154
rect 2620 -1224 2686 -1208
rect 2732 -1154 2798 -1138
rect 2732 -1208 2748 -1154
rect 2782 -1208 2798 -1154
rect 2620 -1274 2692 -1258
rect 2620 -1308 2636 -1274
rect 2670 -1308 2692 -1274
rect 2620 -1324 2692 -1308
rect 2468 -1428 2484 -1374
rect 2518 -1428 2534 -1374
rect 2468 -1444 2534 -1428
rect 2620 -1374 2686 -1358
rect 2620 -1428 2636 -1374
rect 2670 -1428 2686 -1374
rect 2620 -1478 2686 -1428
rect 2732 -1374 2798 -1208
rect 2884 -1154 2950 -1104
rect 2884 -1208 2900 -1154
rect 2934 -1208 2950 -1154
rect 2884 -1224 2950 -1208
rect 2996 -1154 3062 -1138
rect 2996 -1208 3012 -1154
rect 3046 -1208 3062 -1154
rect 2884 -1274 2956 -1258
rect 2884 -1308 2900 -1274
rect 2934 -1308 2956 -1274
rect 2884 -1324 2956 -1308
rect 2732 -1428 2748 -1374
rect 2782 -1428 2798 -1374
rect 2732 -1444 2798 -1428
rect 2884 -1374 2950 -1358
rect 2884 -1428 2900 -1374
rect 2934 -1428 2950 -1374
rect 2884 -1478 2950 -1428
rect 2996 -1374 3062 -1208
rect 3148 -1154 3214 -1104
rect 3148 -1208 3164 -1154
rect 3198 -1208 3214 -1154
rect 3148 -1224 3214 -1208
rect 3260 -1154 3326 -1138
rect 3260 -1208 3276 -1154
rect 3310 -1208 3326 -1154
rect 3148 -1274 3220 -1258
rect 3148 -1308 3164 -1274
rect 3198 -1308 3220 -1274
rect 3148 -1324 3220 -1308
rect 2996 -1428 3012 -1374
rect 3046 -1428 3062 -1374
rect 2996 -1444 3062 -1428
rect 3148 -1374 3214 -1358
rect 3148 -1428 3164 -1374
rect 3198 -1428 3214 -1374
rect 3148 -1478 3214 -1428
rect 3260 -1374 3326 -1208
rect 3412 -1154 3478 -1104
rect 3412 -1208 3428 -1154
rect 3462 -1208 3478 -1154
rect 3412 -1224 3478 -1208
rect 3524 -1154 3590 -1138
rect 3524 -1208 3540 -1154
rect 3574 -1208 3590 -1154
rect 3412 -1274 3484 -1258
rect 3412 -1308 3428 -1274
rect 3462 -1308 3484 -1274
rect 3412 -1324 3484 -1308
rect 3260 -1428 3276 -1374
rect 3310 -1428 3326 -1374
rect 3260 -1444 3326 -1428
rect 3412 -1374 3478 -1358
rect 3412 -1428 3428 -1374
rect 3462 -1428 3478 -1374
rect 3412 -1478 3478 -1428
rect 3524 -1374 3590 -1208
rect 3676 -1154 3742 -1104
rect 3676 -1208 3692 -1154
rect 3726 -1208 3742 -1154
rect 3676 -1224 3742 -1208
rect 3788 -1154 3854 -1138
rect 3788 -1208 3804 -1154
rect 3838 -1208 3854 -1154
rect 3676 -1274 3748 -1258
rect 3676 -1308 3692 -1274
rect 3726 -1308 3748 -1274
rect 3676 -1324 3748 -1308
rect 3524 -1428 3540 -1374
rect 3574 -1428 3590 -1374
rect 3524 -1444 3590 -1428
rect 3676 -1374 3742 -1358
rect 3676 -1428 3692 -1374
rect 3726 -1428 3742 -1374
rect 3676 -1478 3742 -1428
rect 3788 -1374 3854 -1208
rect 3940 -1154 4006 -1104
rect 3940 -1208 3956 -1154
rect 3990 -1208 4006 -1154
rect 3940 -1224 4006 -1208
rect 4052 -1154 4118 -1138
rect 4052 -1208 4068 -1154
rect 4102 -1208 4118 -1154
rect 3940 -1274 4012 -1258
rect 3940 -1308 3956 -1274
rect 3990 -1308 4012 -1274
rect 3940 -1324 4012 -1308
rect 3788 -1428 3804 -1374
rect 3838 -1428 3854 -1374
rect 3788 -1444 3854 -1428
rect 3940 -1374 4006 -1358
rect 3940 -1428 3956 -1374
rect 3990 -1428 4006 -1374
rect 3940 -1478 4006 -1428
rect 4052 -1374 4118 -1208
rect 4052 -1428 4068 -1374
rect 4102 -1428 4118 -1374
rect 4052 -1444 4118 -1428
rect 24 -1498 4170 -1478
rect 24 -1554 72 -1498
rect 4122 -1554 4170 -1498
rect 24 -1574 4170 -1554
rect 24 -1632 120 -1574
rect 24 -2060 46 -1632
rect 100 -1722 120 -1632
rect 226 -1624 292 -1608
rect 226 -1658 242 -1624
rect 276 -1658 292 -1624
rect 226 -1674 292 -1658
rect 358 -1624 424 -1608
rect 358 -1658 374 -1624
rect 408 -1658 424 -1624
rect 358 -1674 424 -1658
rect 490 -1624 556 -1608
rect 490 -1658 506 -1624
rect 540 -1658 556 -1624
rect 490 -1674 556 -1658
rect 622 -1624 688 -1608
rect 622 -1658 638 -1624
rect 672 -1658 688 -1624
rect 622 -1674 688 -1658
rect 754 -1624 820 -1608
rect 754 -1658 770 -1624
rect 804 -1658 820 -1624
rect 754 -1674 820 -1658
rect 886 -1624 952 -1608
rect 886 -1658 902 -1624
rect 936 -1658 952 -1624
rect 886 -1674 952 -1658
rect 1018 -1624 1084 -1608
rect 1018 -1658 1034 -1624
rect 1068 -1658 1084 -1624
rect 1018 -1674 1084 -1658
rect 1150 -1624 1216 -1608
rect 1150 -1658 1166 -1624
rect 1200 -1658 1216 -1624
rect 1150 -1674 1216 -1658
rect 1282 -1624 1348 -1608
rect 1282 -1658 1298 -1624
rect 1332 -1658 1348 -1624
rect 1282 -1674 1348 -1658
rect 1414 -1624 1480 -1608
rect 1414 -1658 1430 -1624
rect 1464 -1658 1480 -1624
rect 1414 -1674 1480 -1658
rect 1546 -1624 1612 -1608
rect 1546 -1658 1562 -1624
rect 1596 -1658 1612 -1624
rect 1546 -1674 1612 -1658
rect 1678 -1624 1744 -1608
rect 1678 -1658 1694 -1624
rect 1728 -1658 1744 -1624
rect 1678 -1674 1744 -1658
rect 1810 -1624 1876 -1608
rect 1810 -1658 1826 -1624
rect 1860 -1658 1876 -1624
rect 1810 -1674 1876 -1658
rect 1942 -1624 2008 -1608
rect 1942 -1658 1958 -1624
rect 1992 -1658 2008 -1624
rect 1942 -1674 2008 -1658
rect 2336 -1624 2402 -1608
rect 2336 -1658 2352 -1624
rect 2386 -1658 2402 -1624
rect 2336 -1674 2402 -1658
rect 2468 -1624 2534 -1608
rect 2468 -1658 2484 -1624
rect 2518 -1658 2534 -1624
rect 2468 -1674 2534 -1658
rect 2600 -1624 2666 -1608
rect 2600 -1658 2616 -1624
rect 2650 -1658 2666 -1624
rect 2600 -1674 2666 -1658
rect 2732 -1624 2798 -1608
rect 2732 -1658 2748 -1624
rect 2782 -1658 2798 -1624
rect 2732 -1674 2798 -1658
rect 2864 -1624 2930 -1608
rect 2864 -1658 2880 -1624
rect 2914 -1658 2930 -1624
rect 2864 -1674 2930 -1658
rect 2996 -1624 3062 -1608
rect 2996 -1658 3012 -1624
rect 3046 -1658 3062 -1624
rect 2996 -1674 3062 -1658
rect 3128 -1624 3194 -1608
rect 3128 -1658 3144 -1624
rect 3178 -1658 3194 -1624
rect 3128 -1674 3194 -1658
rect 3260 -1624 3326 -1608
rect 3260 -1658 3276 -1624
rect 3310 -1658 3326 -1624
rect 3260 -1674 3326 -1658
rect 3392 -1624 3458 -1608
rect 3392 -1658 3408 -1624
rect 3442 -1658 3458 -1624
rect 3392 -1674 3458 -1658
rect 3524 -1624 3590 -1608
rect 3524 -1658 3540 -1624
rect 3574 -1658 3590 -1624
rect 3524 -1674 3590 -1658
rect 3656 -1624 3722 -1608
rect 3656 -1658 3672 -1624
rect 3706 -1658 3722 -1624
rect 3656 -1674 3722 -1658
rect 3788 -1624 3854 -1608
rect 3788 -1658 3804 -1624
rect 3838 -1658 3854 -1624
rect 3788 -1674 3854 -1658
rect 3920 -1624 3986 -1608
rect 3920 -1658 3936 -1624
rect 3970 -1658 3986 -1624
rect 3920 -1674 3986 -1658
rect 4052 -1624 4118 -1608
rect 4052 -1658 4068 -1624
rect 4102 -1658 4118 -1624
rect 4052 -1674 4118 -1658
rect 100 -1738 358 -1722
rect 100 -1792 176 -1738
rect 210 -1792 308 -1738
rect 342 -1792 358 -1738
rect 100 -1808 358 -1792
rect 424 -1738 622 -1722
rect 424 -1792 440 -1738
rect 474 -1792 572 -1738
rect 606 -1792 622 -1738
rect 424 -1808 622 -1792
rect 688 -1738 886 -1722
rect 688 -1792 704 -1738
rect 738 -1792 836 -1738
rect 870 -1792 886 -1738
rect 688 -1808 886 -1792
rect 952 -1738 1150 -1722
rect 952 -1792 968 -1738
rect 1002 -1792 1100 -1738
rect 1134 -1792 1150 -1738
rect 952 -1808 1150 -1792
rect 1216 -1738 1414 -1722
rect 1216 -1792 1232 -1738
rect 1266 -1792 1364 -1738
rect 1398 -1792 1414 -1738
rect 1216 -1808 1414 -1792
rect 1480 -1738 1678 -1722
rect 1480 -1792 1496 -1738
rect 1530 -1792 1628 -1738
rect 1662 -1792 1678 -1738
rect 1480 -1808 1678 -1792
rect 1744 -1738 1942 -1722
rect 1744 -1792 1760 -1738
rect 1794 -1792 1892 -1738
rect 1926 -1792 1942 -1738
rect 1744 -1808 1942 -1792
rect 2008 -1738 2336 -1722
rect 2008 -1792 2024 -1738
rect 2058 -1792 2286 -1738
rect 2320 -1792 2336 -1738
rect 2008 -1808 2336 -1792
rect 2402 -1738 2468 -1722
rect 2402 -1792 2418 -1738
rect 2452 -1792 2468 -1738
rect 100 -1864 120 -1808
rect 100 -1880 358 -1864
rect 100 -1934 176 -1880
rect 210 -1934 308 -1880
rect 342 -1934 358 -1880
rect 100 -1950 358 -1934
rect 424 -1880 622 -1864
rect 424 -1934 440 -1880
rect 474 -1934 572 -1880
rect 606 -1934 622 -1880
rect 424 -1950 622 -1934
rect 688 -1880 886 -1864
rect 688 -1934 704 -1880
rect 738 -1934 836 -1880
rect 870 -1934 886 -1880
rect 688 -1950 886 -1934
rect 952 -1880 1150 -1864
rect 952 -1934 968 -1880
rect 1002 -1934 1100 -1880
rect 1134 -1934 1150 -1880
rect 952 -1950 1150 -1934
rect 1216 -1880 1414 -1864
rect 1216 -1934 1232 -1880
rect 1266 -1934 1364 -1880
rect 1398 -1934 1414 -1880
rect 1216 -1950 1414 -1934
rect 1480 -1880 1678 -1864
rect 1480 -1934 1496 -1880
rect 1530 -1934 1628 -1880
rect 1662 -1934 1678 -1880
rect 1480 -1950 1678 -1934
rect 1744 -1880 1810 -1864
rect 1744 -1934 1760 -1880
rect 1794 -1934 1810 -1880
rect 1744 -1950 1810 -1934
rect 1876 -1880 2336 -1864
rect 1876 -1934 1892 -1880
rect 1926 -1934 2024 -1880
rect 2058 -1934 2286 -1880
rect 2320 -1934 2336 -1880
rect 1876 -1950 2336 -1934
rect 2402 -1880 2468 -1792
rect 2534 -1738 2600 -1722
rect 2534 -1792 2550 -1738
rect 2584 -1792 2600 -1738
rect 2534 -1808 2600 -1792
rect 2666 -1738 2732 -1722
rect 2666 -1792 2682 -1738
rect 2716 -1792 2732 -1738
rect 2402 -1934 2418 -1880
rect 2452 -1934 2468 -1880
rect 100 -2060 120 -1950
rect 24 -2116 120 -2060
rect 2402 -2124 2468 -1934
rect 2534 -1880 2600 -1864
rect 2534 -1934 2550 -1880
rect 2584 -1934 2600 -1880
rect 2534 -1950 2600 -1934
rect 2666 -1880 2732 -1792
rect 2798 -1738 2864 -1722
rect 2798 -1792 2814 -1738
rect 2848 -1792 2864 -1738
rect 2798 -1808 2864 -1792
rect 2930 -1738 2996 -1722
rect 2930 -1792 2946 -1738
rect 2980 -1792 2996 -1738
rect 2666 -1934 2682 -1880
rect 2716 -1934 2732 -1880
rect 2666 -2124 2732 -1934
rect 2798 -1880 2864 -1864
rect 2798 -1934 2814 -1880
rect 2848 -1934 2864 -1880
rect 2798 -1950 2864 -1934
rect 2930 -1880 2996 -1792
rect 3062 -1738 3128 -1722
rect 3062 -1792 3078 -1738
rect 3112 -1792 3128 -1738
rect 3062 -1808 3128 -1792
rect 3194 -1738 3260 -1722
rect 3194 -1792 3210 -1738
rect 3244 -1792 3260 -1738
rect 2930 -1934 2946 -1880
rect 2980 -1934 2996 -1880
rect 2930 -2124 2996 -1934
rect 3062 -1880 3128 -1864
rect 3062 -1934 3078 -1880
rect 3112 -1934 3128 -1880
rect 3062 -1950 3128 -1934
rect 3194 -1880 3260 -1792
rect 3326 -1738 3392 -1722
rect 3326 -1792 3342 -1738
rect 3376 -1792 3392 -1738
rect 3326 -1808 3392 -1792
rect 3458 -1738 3524 -1722
rect 3458 -1792 3474 -1738
rect 3508 -1792 3524 -1738
rect 3194 -1934 3210 -1880
rect 3244 -1934 3260 -1880
rect 3194 -2124 3260 -1934
rect 3326 -1880 3392 -1864
rect 3326 -1934 3342 -1880
rect 3376 -1934 3392 -1880
rect 3326 -1950 3392 -1934
rect 3458 -1880 3524 -1792
rect 3590 -1738 3656 -1722
rect 3590 -1792 3606 -1738
rect 3640 -1792 3656 -1738
rect 3590 -1808 3656 -1792
rect 3722 -1738 3788 -1722
rect 3722 -1792 3738 -1738
rect 3772 -1792 3788 -1738
rect 3458 -1934 3474 -1880
rect 3508 -1934 3524 -1880
rect 3458 -2124 3524 -1934
rect 3590 -1880 3656 -1864
rect 3590 -1934 3606 -1880
rect 3640 -1934 3656 -1880
rect 3590 -1950 3656 -1934
rect 3722 -1880 3788 -1792
rect 3854 -1738 3920 -1722
rect 3854 -1792 3870 -1738
rect 3904 -1792 3920 -1738
rect 3854 -1808 3920 -1792
rect 3986 -1738 4052 -1722
rect 3986 -1792 4002 -1738
rect 4036 -1792 4052 -1738
rect 3722 -1934 3738 -1880
rect 3772 -1934 3788 -1880
rect 3722 -2124 3788 -1934
rect 3854 -1880 3920 -1864
rect 3854 -1934 3870 -1880
rect 3904 -1934 3920 -1880
rect 3854 -1950 3920 -1934
rect 3986 -1880 4052 -1792
rect 3986 -1934 4002 -1880
rect 4036 -1934 4052 -1880
rect 3986 -2124 4052 -1934
rect 4204 -2124 4294 -1104
rect 2138 -2144 4294 -2124
rect 2138 -2200 2186 -2144
rect 4090 -2200 4294 -2144
rect 2138 -2220 4294 -2200
<< viali >>
rect 354 -1308 388 -1274
rect 242 -1428 276 -1374
rect 618 -1308 652 -1274
rect 506 -1428 540 -1374
rect 882 -1308 916 -1274
rect 770 -1428 804 -1374
rect 1146 -1308 1180 -1274
rect 1034 -1428 1068 -1374
rect 1410 -1308 1444 -1274
rect 1298 -1428 1332 -1374
rect 1674 -1308 1708 -1274
rect 1562 -1428 1596 -1374
rect 1938 -1308 1972 -1274
rect 2372 -1308 2406 -1274
rect 1826 -1428 1860 -1374
rect 2636 -1308 2670 -1274
rect 2484 -1428 2518 -1374
rect 2900 -1308 2934 -1274
rect 2748 -1428 2782 -1374
rect 3164 -1308 3198 -1274
rect 3012 -1428 3046 -1374
rect 3428 -1308 3462 -1274
rect 3276 -1428 3310 -1374
rect 3692 -1308 3726 -1274
rect 3540 -1428 3574 -1374
rect 3956 -1308 3990 -1274
rect 3804 -1428 3838 -1374
rect 4068 -1428 4102 -1374
rect 242 -1658 276 -1624
rect 374 -1658 408 -1624
rect 506 -1658 540 -1624
rect 638 -1658 672 -1624
rect 770 -1658 804 -1624
rect 902 -1658 936 -1624
rect 1034 -1658 1068 -1624
rect 1166 -1658 1200 -1624
rect 1298 -1658 1332 -1624
rect 1430 -1658 1464 -1624
rect 1562 -1658 1596 -1624
rect 1694 -1658 1728 -1624
rect 1826 -1658 1860 -1624
rect 1958 -1658 1992 -1624
rect 2352 -1658 2386 -1624
rect 2484 -1658 2518 -1624
rect 2616 -1658 2650 -1624
rect 2748 -1658 2782 -1624
rect 2880 -1658 2914 -1624
rect 3012 -1658 3046 -1624
rect 3144 -1658 3178 -1624
rect 3276 -1658 3310 -1624
rect 3408 -1658 3442 -1624
rect 3540 -1658 3574 -1624
rect 3672 -1658 3706 -1624
rect 3804 -1658 3838 -1624
rect 3936 -1658 3970 -1624
rect 4068 -1658 4102 -1624
rect 2286 -1792 2320 -1738
rect 2286 -1934 2320 -1880
rect 2550 -1792 2584 -1738
rect 2550 -1934 2584 -1880
rect 2814 -1792 2848 -1738
rect 2814 -1934 2848 -1880
rect 3078 -1792 3112 -1738
rect 3078 -1934 3112 -1880
rect 3342 -1792 3376 -1738
rect 3342 -1934 3376 -1880
rect 3606 -1792 3640 -1738
rect 3606 -1934 3640 -1880
rect 3870 -1792 3904 -1738
rect 3870 -1934 3904 -1880
<< metal1 >>
rect 353 -700 3991 -694
rect 353 -754 434 -700
rect 498 -754 3991 -700
rect 353 -760 3991 -754
rect 353 -1258 419 -760
rect 619 -794 3725 -788
rect 619 -848 708 -794
rect 772 -848 3725 -794
rect 619 -854 3725 -848
rect 619 -1258 685 -854
rect 891 -888 3457 -882
rect 891 -942 964 -888
rect 1028 -942 3457 -888
rect 891 -948 3457 -942
rect 891 -1258 957 -948
rect 1150 -982 3194 -976
rect 1150 -1036 1226 -982
rect 1290 -1036 3194 -982
rect 1150 -1042 3194 -1036
rect 1150 -1258 1216 -1042
rect 1414 -1076 2932 -1070
rect 1414 -1130 1488 -1076
rect 1552 -1130 2932 -1076
rect 1414 -1136 2932 -1130
rect 1414 -1258 1480 -1136
rect 1678 -1170 2666 -1164
rect 1678 -1224 1752 -1170
rect 1816 -1224 2666 -1170
rect 1678 -1230 2666 -1224
rect 1678 -1258 1744 -1230
rect 2600 -1258 2666 -1230
rect 2864 -1258 2932 -1136
rect 3126 -1258 3194 -1042
rect 3391 -1258 3457 -948
rect 3659 -1258 3725 -854
rect 3925 -1258 3991 -760
rect 338 -1274 424 -1258
rect 338 -1308 354 -1274
rect 388 -1308 424 -1274
rect 338 -1324 424 -1308
rect 602 -1274 688 -1258
rect 602 -1308 618 -1274
rect 652 -1308 688 -1274
rect 602 -1324 688 -1308
rect 866 -1274 957 -1258
rect 866 -1308 882 -1274
rect 916 -1308 957 -1274
rect 866 -1321 957 -1308
rect 1130 -1274 1216 -1258
rect 1130 -1308 1146 -1274
rect 1180 -1308 1216 -1274
rect 866 -1324 952 -1321
rect 1130 -1324 1216 -1308
rect 1394 -1274 1480 -1258
rect 1394 -1308 1410 -1274
rect 1444 -1308 1480 -1274
rect 1394 -1324 1480 -1308
rect 1658 -1274 1744 -1258
rect 1658 -1308 1674 -1274
rect 1708 -1308 1744 -1274
rect 1658 -1324 1744 -1308
rect 1922 -1264 2422 -1258
rect 1922 -1274 2030 -1264
rect 1922 -1308 1938 -1274
rect 1972 -1308 2030 -1274
rect 1922 -1318 2030 -1308
rect 2094 -1274 2422 -1264
rect 2094 -1308 2372 -1274
rect 2406 -1308 2422 -1274
rect 2094 -1318 2422 -1308
rect 1922 -1324 2422 -1318
rect 2600 -1274 2686 -1258
rect 2600 -1308 2636 -1274
rect 2670 -1308 2686 -1274
rect 2600 -1324 2686 -1308
rect 2864 -1274 2950 -1258
rect 2864 -1308 2900 -1274
rect 2934 -1308 2950 -1274
rect 3126 -1274 3214 -1258
rect 3126 -1292 3164 -1274
rect 2864 -1324 2950 -1308
rect 3128 -1308 3164 -1292
rect 3198 -1308 3214 -1274
rect 3128 -1324 3214 -1308
rect 3391 -1274 3478 -1258
rect 3391 -1308 3428 -1274
rect 3462 -1308 3478 -1274
rect 3391 -1313 3478 -1308
rect 3392 -1324 3478 -1313
rect 3656 -1274 3742 -1258
rect 3656 -1308 3692 -1274
rect 3726 -1308 3742 -1274
rect 3656 -1324 3742 -1308
rect 3920 -1274 4006 -1258
rect 3920 -1308 3956 -1274
rect 3990 -1308 4006 -1274
rect 3920 -1324 4006 -1308
rect 353 -1327 424 -1324
rect 226 -1374 292 -1358
rect 226 -1428 242 -1374
rect 276 -1428 292 -1374
rect 226 -1624 292 -1428
rect 226 -1658 242 -1624
rect 276 -1658 292 -1624
rect 226 -1674 292 -1658
rect 358 -1624 424 -1327
rect 358 -1658 374 -1624
rect 408 -1658 424 -1624
rect 358 -1674 424 -1658
rect 490 -1374 556 -1358
rect 490 -1428 506 -1374
rect 540 -1428 556 -1374
rect 490 -1624 556 -1428
rect 490 -1658 506 -1624
rect 540 -1658 556 -1624
rect 490 -1674 556 -1658
rect 622 -1624 688 -1324
rect 622 -1658 638 -1624
rect 672 -1658 688 -1624
rect 622 -1674 688 -1658
rect 754 -1374 820 -1358
rect 754 -1428 770 -1374
rect 804 -1428 820 -1374
rect 754 -1624 820 -1428
rect 754 -1658 770 -1624
rect 804 -1658 820 -1624
rect 754 -1674 820 -1658
rect 886 -1624 952 -1324
rect 886 -1658 902 -1624
rect 936 -1658 952 -1624
rect 886 -1674 952 -1658
rect 1018 -1374 1084 -1358
rect 1018 -1428 1034 -1374
rect 1068 -1428 1084 -1374
rect 1018 -1624 1084 -1428
rect 1018 -1658 1034 -1624
rect 1068 -1658 1084 -1624
rect 1018 -1674 1084 -1658
rect 1150 -1624 1216 -1324
rect 1150 -1658 1166 -1624
rect 1200 -1658 1216 -1624
rect 1150 -1674 1216 -1658
rect 1282 -1374 1348 -1358
rect 1282 -1428 1298 -1374
rect 1332 -1428 1348 -1374
rect 1282 -1624 1348 -1428
rect 1282 -1658 1298 -1624
rect 1332 -1658 1348 -1624
rect 1282 -1674 1348 -1658
rect 1414 -1624 1480 -1324
rect 1414 -1658 1430 -1624
rect 1464 -1658 1480 -1624
rect 1414 -1674 1480 -1658
rect 1546 -1374 1612 -1358
rect 1546 -1428 1562 -1374
rect 1596 -1428 1612 -1374
rect 1546 -1624 1612 -1428
rect 1546 -1658 1562 -1624
rect 1596 -1658 1612 -1624
rect 1546 -1674 1612 -1658
rect 1678 -1624 1744 -1324
rect 1678 -1658 1694 -1624
rect 1728 -1658 1744 -1624
rect 1678 -1674 1744 -1658
rect 1810 -1374 1876 -1358
rect 1810 -1428 1826 -1374
rect 1860 -1428 1876 -1374
rect 1810 -1624 1876 -1428
rect 1810 -1658 1826 -1624
rect 1860 -1658 1876 -1624
rect 1810 -1674 1876 -1658
rect 1942 -1624 2008 -1324
rect 1942 -1658 1958 -1624
rect 1992 -1658 2008 -1624
rect 1942 -1674 2008 -1658
rect 2336 -1624 2402 -1324
rect 2336 -1658 2352 -1624
rect 2386 -1658 2402 -1624
rect 2336 -1674 2402 -1658
rect 2468 -1374 2534 -1358
rect 2468 -1428 2484 -1374
rect 2518 -1428 2534 -1374
rect 2468 -1624 2534 -1428
rect 2468 -1658 2484 -1624
rect 2518 -1658 2534 -1624
rect 2468 -1674 2534 -1658
rect 2600 -1624 2666 -1324
rect 2600 -1658 2616 -1624
rect 2650 -1658 2666 -1624
rect 2600 -1674 2666 -1658
rect 2732 -1374 2798 -1358
rect 2732 -1428 2748 -1374
rect 2782 -1428 2798 -1374
rect 2732 -1624 2798 -1428
rect 2732 -1658 2748 -1624
rect 2782 -1658 2798 -1624
rect 2732 -1674 2798 -1658
rect 2864 -1624 2930 -1324
rect 2864 -1658 2880 -1624
rect 2914 -1658 2930 -1624
rect 2864 -1674 2930 -1658
rect 2996 -1374 3062 -1358
rect 2996 -1428 3012 -1374
rect 3046 -1428 3062 -1374
rect 2996 -1624 3062 -1428
rect 2996 -1658 3012 -1624
rect 3046 -1658 3062 -1624
rect 2996 -1674 3062 -1658
rect 3128 -1624 3194 -1324
rect 3128 -1658 3144 -1624
rect 3178 -1658 3194 -1624
rect 3128 -1674 3194 -1658
rect 3260 -1374 3326 -1358
rect 3260 -1428 3276 -1374
rect 3310 -1428 3326 -1374
rect 3260 -1624 3326 -1428
rect 3260 -1658 3276 -1624
rect 3310 -1658 3326 -1624
rect 3260 -1674 3326 -1658
rect 3392 -1624 3458 -1324
rect 3392 -1658 3408 -1624
rect 3442 -1658 3458 -1624
rect 3392 -1674 3458 -1658
rect 3524 -1374 3590 -1358
rect 3524 -1428 3540 -1374
rect 3574 -1428 3590 -1374
rect 3524 -1624 3590 -1428
rect 3524 -1658 3540 -1624
rect 3574 -1658 3590 -1624
rect 3524 -1674 3590 -1658
rect 3656 -1624 3722 -1324
rect 3920 -1327 3991 -1324
rect 3656 -1658 3672 -1624
rect 3706 -1658 3722 -1624
rect 3656 -1674 3722 -1658
rect 3788 -1374 3854 -1358
rect 3788 -1428 3804 -1374
rect 3838 -1428 3854 -1374
rect 3788 -1624 3854 -1428
rect 3788 -1658 3804 -1624
rect 3838 -1658 3854 -1624
rect 3788 -1674 3854 -1658
rect 3920 -1624 3986 -1327
rect 3920 -1658 3936 -1624
rect 3970 -1658 3986 -1624
rect 3920 -1674 3986 -1658
rect 4052 -1374 4118 -1358
rect 4052 -1428 4068 -1374
rect 4102 -1428 4118 -1374
rect 4052 -1624 4118 -1428
rect 4052 -1658 4068 -1624
rect 4102 -1658 4118 -1624
rect 4052 -1674 4118 -1658
rect 2270 -1738 4294 -1722
rect 2270 -1792 2286 -1738
rect 2320 -1792 2550 -1738
rect 2584 -1792 2814 -1738
rect 2848 -1792 3078 -1738
rect 3112 -1792 3342 -1738
rect 3376 -1792 3606 -1738
rect 3640 -1792 3870 -1738
rect 3904 -1792 4294 -1738
rect 2270 -1808 4294 -1792
rect 2270 -1880 4294 -1864
rect 2270 -1934 2286 -1880
rect 2320 -1934 2550 -1880
rect 2584 -1934 2814 -1880
rect 2848 -1934 3078 -1880
rect 3112 -1934 3342 -1880
rect 3376 -1934 3606 -1880
rect 3640 -1934 3870 -1880
rect 3904 -1934 4294 -1880
rect 2270 -1950 4294 -1934
<< via1 >>
rect 434 -754 498 -700
rect 708 -848 772 -794
rect 964 -942 1028 -888
rect 1226 -1036 1290 -982
rect 1488 -1130 1552 -1076
rect 1752 -1224 1816 -1170
rect 2030 -1318 2094 -1264
<< metal2 >>
rect 428 -700 504 -694
rect 428 -754 434 -700
rect 498 -754 504 -700
rect 428 -760 504 -754
rect 702 -794 778 -788
rect 702 -848 708 -794
rect 772 -848 778 -794
rect 702 -854 778 -848
rect 958 -888 1034 -882
rect 958 -942 964 -888
rect 1028 -942 1034 -888
rect 958 -948 1034 -942
rect 1220 -982 1296 -976
rect 1220 -1036 1226 -982
rect 1290 -1036 1296 -982
rect 1220 -1042 1296 -1036
rect 1482 -1076 1558 -1070
rect 1482 -1130 1488 -1076
rect 1552 -1130 1558 -1076
rect 1482 -1136 1558 -1130
rect 1746 -1170 1822 -1164
rect 1746 -1224 1752 -1170
rect 1816 -1224 1822 -1170
rect 1746 -1230 1822 -1224
rect 2024 -1264 2100 -1258
rect 2024 -1318 2030 -1264
rect 2094 -1318 2100 -1264
rect 2024 -1324 2100 -1318
<< labels >>
flabel locali 4204 -1644 4294 -1104 0 FreeSerif 160 0 0 0 GND!
port 50 nsew
flabel locali 24 -2116 120 -1576 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel metal1 4204 -1808 4294 -1722 0 FreeSerif 160 0 0 0 word0
port 36 nsew
flabel metal1 4204 -1950 4294 -1864 0 FreeSerif 160 0 0 0 word1
port 65 nsew
flabel metal2 428 -760 504 -694 0 FreeSerif 160 0 0 0 A6
port 14 nsew
flabel metal2 702 -854 778 -788 0 FreeSerif 160 0 0 0 A5
port 13 nsew
flabel metal2 958 -948 1034 -882 0 FreeSerif 160 0 0 0 A4
port 12 nsew
flabel metal2 1220 -1042 1296 -976 0 FreeSerif 160 0 0 0 A3
port 11 nsew
flabel metal2 1482 -1136 1558 -1070 0 FreeSerif 160 0 0 0 A2
port 10 nsew
flabel metal2 1746 -1230 1822 -1164 0 FreeSerif 160 0 0 0 A1
port 9 nsew
flabel metal2 2024 -1324 2100 -1258 0 FreeSerif 160 0 0 0 A0
port 8 nsew
<< end >>
