magic
tech sky130A
magscale 1 2
timestamp 1745485683
<< locali >>
rect -314 864 12226 960
rect 2685 693 2739 747
rect 5923 693 5977 747
rect 9161 693 9215 747
rect 3104 498 3170 692
rect 1010 374 1062 426
rect 4248 374 4300 426
rect 6342 474 6408 668
rect 9580 488 9646 682
rect 7486 374 7538 426
rect 10724 374 10776 426
rect 11902 370 11968 436
rect 1738 306 1792 358
rect 2788 304 3068 368
rect 3104 295 3343 361
rect 4976 306 5030 358
rect 6026 304 6306 368
rect 6342 291 6593 357
rect 8214 306 8268 358
rect 9264 304 9544 368
rect 9580 293 9847 359
rect 11452 306 11506 358
rect -314 0 12226 96
<< viali >>
rect 88 625 142 679
rect -130 414 -90 454
rect 2689 423 2743 477
rect 2202 384 2240 422
rect 5929 423 5983 477
rect 9165 427 9219 481
rect 5440 384 5478 422
rect 8678 384 8716 422
rect -231 299 -177 353
rect 2581 301 2635 355
rect 5819 301 5873 355
rect 9057 301 9111 355
<< metal1 >>
rect 82 679 148 691
rect 82 625 88 679
rect 142 625 148 679
rect 82 529 148 625
rect 407 531 413 597
rect 479 531 485 597
rect 2549 523 2555 589
rect 2621 523 2627 589
rect 3645 531 3651 597
rect 3717 531 3723 597
rect 2555 483 2621 523
rect 5804 521 5810 587
rect 5876 521 5882 587
rect 6883 531 6889 597
rect 6955 531 6961 597
rect 9040 521 9046 587
rect 9112 521 9118 587
rect 10121 531 10199 597
rect 5810 483 5876 521
rect 9046 487 9112 521
rect 2555 477 2755 483
rect -136 460 -84 466
rect -136 402 -84 408
rect 2188 422 2457 436
rect 2188 384 2202 422
rect 2240 384 2457 422
rect 2555 423 2689 477
rect 2743 423 2755 477
rect 5810 477 5995 483
rect 2555 417 2755 423
rect 2188 370 2457 384
rect 5426 422 5695 436
rect 5426 384 5440 422
rect 5478 384 5695 422
rect 5810 423 5929 477
rect 5983 423 5995 477
rect 9046 481 9231 487
rect 5810 417 5995 423
rect 5426 370 5695 384
rect 8664 422 8933 436
rect 8664 384 8678 422
rect 8716 384 8933 422
rect 9046 427 9165 481
rect 9219 427 9231 481
rect 9046 421 9231 427
rect 8664 370 8933 384
rect -237 359 -171 365
rect 2391 361 2457 370
rect 5629 361 5695 370
rect 8867 361 8933 370
rect 2391 355 2647 361
rect 2391 301 2581 355
rect 2635 301 2647 355
rect 5629 355 5885 361
rect 2391 295 2647 301
rect 5629 301 5819 355
rect 5873 301 5885 355
rect 8867 355 9123 361
rect 5629 295 5885 301
rect 8867 301 9057 355
rect 9111 301 9123 355
rect 8867 295 9123 301
rect -237 287 -171 293
<< via1 >>
rect 413 531 479 597
rect 2555 523 2621 589
rect 3651 531 3717 597
rect 5810 521 5876 587
rect 6889 531 6955 597
rect 9046 521 9112 587
rect -136 454 -84 460
rect -136 414 -130 454
rect -130 414 -90 454
rect -90 414 -84 454
rect -136 408 -84 414
rect 1010 374 1062 426
rect 4248 374 4300 426
rect 7486 374 7538 426
rect 10724 374 10776 426
rect -237 353 -171 359
rect -237 299 -231 353
rect -231 299 -177 353
rect -177 299 -171 353
rect 1738 306 1792 358
rect -237 293 -171 299
rect 4976 306 5030 358
rect 8214 306 8268 358
rect 11452 306 11506 358
<< metal2 >>
rect 412 687 2622 753
rect 3650 687 5876 753
rect 6888 687 9112 753
rect 413 597 479 687
rect 413 525 479 531
rect 2555 589 2621 687
rect 3651 597 3717 687
rect 3651 525 3717 531
rect 5810 587 5876 687
rect 2555 517 2621 523
rect 6889 597 6955 687
rect 6889 525 6955 531
rect 9046 587 9112 687
rect 5810 515 5876 521
rect 9046 515 9112 521
rect -142 408 -136 460
rect -84 458 -78 460
rect 1018 458 3340 468
rect 7494 458 9800 460
rect -84 410 434 458
rect 1018 432 3672 458
rect 6484 448 6910 458
rect 4252 432 6910 448
rect 7494 432 10148 458
rect -84 408 -78 410
rect 386 374 434 410
rect 1004 426 3672 432
rect 1004 374 1010 426
rect 1062 420 3672 426
rect 1062 374 1070 420
rect 3246 410 3672 420
rect -236 359 -172 362
rect -243 293 -237 359
rect -171 293 5 359
rect 386 326 1070 374
rect 3624 374 3672 410
rect 4242 426 6910 432
rect 4242 374 4248 426
rect 4300 410 6910 426
rect 4300 400 6568 410
rect 4300 374 4308 400
rect 1730 358 1796 366
rect -236 288 -172 293
rect -61 261 5 293
rect 1730 306 1738 358
rect 1792 306 1796 358
rect 3624 326 4308 374
rect 6862 374 6910 410
rect 7480 426 10148 432
rect 7480 374 7486 426
rect 7538 412 10148 426
rect 7538 374 7546 412
rect 9722 410 10148 412
rect 4968 358 5034 366
rect 1730 261 1796 306
rect 4968 306 4976 358
rect 5030 306 5034 358
rect 6862 326 7546 374
rect 10100 374 10148 410
rect 10718 426 10784 432
rect 10718 374 10724 426
rect 10776 374 10784 426
rect 8206 358 8272 366
rect 4968 261 5034 306
rect 8206 306 8214 358
rect 8268 306 8272 358
rect 10100 326 10784 374
rect 11444 358 11510 366
rect 8206 261 8272 306
rect 11444 306 11452 358
rect 11506 306 11510 358
rect 11444 261 11510 306
rect -61 195 11510 261
use inv  inv_1 ~/magic/library/mag
timestamp 1738780557
transform 1 0 -314 0 1 0
box -4 0 322 976
use inv  inv_2
timestamp 1738780557
transform 1 0 2924 0 1 0
box -4 0 322 976
use inv  inv_3
timestamp 1738780557
transform 1 0 6162 0 1 0
box -4 0 322 976
use inv  inv_4
timestamp 1738780557
transform 1 0 9400 0 1 0
box -4 0 322 976
use nand  nand_0 ~/magic/library/mag
timestamp 1739944168
transform 1 0 8974 0 1 0
box -4 0 430 976
use nand  nand_1
timestamp 1739944168
transform 1 0 2498 0 1 0
box -4 0 430 976
use nand  nand_2
timestamp 1739944168
transform 1 0 5736 0 1 0
box -4 0 430 976
use tff  tff_0
timestamp 1745480928
transform 1 0 6776 0 1 0
box -300 0 2212 976
use tff  tff_1
timestamp 1745480928
transform 1 0 300 0 1 0
box -300 0 2212 976
use tff  tff_2
timestamp 1745480928
transform 1 0 3538 0 1 0
box -300 0 2212 976
use tff  tff_3
timestamp 1745480928
transform 1 0 10014 0 1 0
box -300 0 2212 976
<< labels >>
flabel locali -314 864 12226 960 0 FreeSerif 160 0 0 0 VDD!
flabel locali -314 0 12226 96 0 FreeSerif 160 0 0 0 GND!
flabel metal2 -236 288 -172 362 0 FreeSerif 160 0 0 0 CLK
port 2 nsew
flabel metal1 2391 296 2502 360 0 FreeSerif 160 0 0 0 Q0
port 5 nsew
flabel metal1 5630 296 5774 360 0 FreeSerif 160 0 0 0 Q1
port 9 nsew
flabel metal1 8870 296 9008 360 0 FreeSerif 160 0 0 0 Q2
port 13 nsew
flabel locali 11902 370 11968 436 0 FreeSerif 160 0 0 0 Q3
port 16 nsew
<< end >>
