magic
tech sky130A
magscale 1 2
timestamp 1744932088
<< nwell >>
rect -54 -17710 1946 -17350
<< nmos >>
rect 978 -17986 1080 -17952
rect 1476 -17986 1578 -17952
rect 1476 -18128 1578 -18094
<< pmos >>
rect -18 -17602 84 -17568
rect 314 -17602 416 -17568
rect 480 -17602 582 -17568
rect 812 -17602 914 -17568
rect 978 -17602 1080 -17568
rect 1310 -17602 1412 -17568
rect 1476 -17602 1578 -17568
rect 1808 -17602 1910 -17568
<< ndiff >>
rect 978 -17880 1080 -17864
rect 978 -17914 1012 -17880
rect 1046 -17914 1080 -17880
rect 978 -17952 1080 -17914
rect 1476 -17880 1578 -17864
rect 1476 -17914 1510 -17880
rect 1544 -17914 1578 -17880
rect 1476 -17952 1578 -17914
rect 978 -18006 1080 -17986
rect 1476 -18006 1578 -17986
rect 978 -18022 1228 -18006
rect 978 -18056 1178 -18022
rect 1212 -18056 1228 -18022
rect 978 -18072 1228 -18056
rect 1476 -18022 1726 -18006
rect 1476 -18056 1676 -18022
rect 1710 -18056 1726 -18022
rect 1476 -18072 1726 -18056
rect 1476 -18094 1578 -18072
rect 1476 -18164 1578 -18128
rect 1476 -18198 1510 -18164
rect 1544 -18198 1578 -18164
rect 1476 -18214 1578 -18198
<< pdiff >>
rect -18 -17512 84 -17496
rect -18 -17546 -2 -17512
rect 66 -17546 84 -17512
rect -18 -17568 84 -17546
rect 314 -17512 416 -17496
rect 314 -17546 330 -17512
rect 398 -17546 416 -17512
rect 314 -17568 416 -17546
rect 480 -17512 582 -17496
rect 480 -17546 496 -17512
rect 564 -17546 582 -17512
rect 480 -17568 582 -17546
rect 812 -17512 914 -17496
rect 812 -17546 828 -17512
rect 896 -17546 914 -17512
rect 812 -17568 914 -17546
rect 978 -17512 1080 -17496
rect 978 -17546 994 -17512
rect 1062 -17546 1080 -17512
rect 978 -17568 1080 -17546
rect 1310 -17512 1412 -17496
rect 1310 -17546 1326 -17512
rect 1394 -17546 1412 -17512
rect 1310 -17568 1412 -17546
rect 1476 -17512 1578 -17496
rect 1476 -17546 1492 -17512
rect 1560 -17546 1578 -17512
rect 1476 -17568 1578 -17546
rect 1808 -17512 1910 -17496
rect 1808 -17546 1824 -17512
rect 1892 -17546 1910 -17512
rect 1808 -17568 1910 -17546
rect -18 -17624 84 -17602
rect -18 -17658 16 -17624
rect 50 -17658 84 -17624
rect -18 -17674 84 -17658
rect 314 -17624 416 -17602
rect 314 -17658 348 -17624
rect 382 -17658 416 -17624
rect 314 -17674 416 -17658
rect 480 -17624 582 -17602
rect 480 -17658 514 -17624
rect 548 -17658 582 -17624
rect 480 -17674 582 -17658
rect 812 -17624 914 -17602
rect 812 -17658 846 -17624
rect 880 -17658 914 -17624
rect 812 -17674 914 -17658
rect 978 -17624 1080 -17602
rect 978 -17658 1012 -17624
rect 1046 -17658 1080 -17624
rect 978 -17674 1080 -17658
rect 1310 -17624 1412 -17602
rect 1310 -17658 1344 -17624
rect 1378 -17658 1412 -17624
rect 1310 -17674 1412 -17658
rect 1476 -17624 1578 -17602
rect 1476 -17658 1510 -17624
rect 1544 -17658 1578 -17624
rect 1476 -17674 1578 -17658
rect 1808 -17624 1910 -17602
rect 1808 -17658 1842 -17624
rect 1876 -17658 1910 -17624
rect 1808 -17674 1910 -17658
<< ndiffc >>
rect 1012 -17914 1046 -17880
rect 1510 -17914 1544 -17880
rect 1178 -18056 1212 -18022
rect 1676 -18056 1710 -18022
rect 1510 -18198 1544 -18164
<< pdiffc >>
rect -2 -17546 66 -17512
rect 330 -17546 398 -17512
rect 496 -17546 564 -17512
rect 828 -17546 896 -17512
rect 994 -17546 1062 -17512
rect 1326 -17546 1394 -17512
rect 1492 -17546 1560 -17512
rect 1824 -17546 1892 -17512
rect 16 -17658 50 -17624
rect 348 -17658 382 -17624
rect 514 -17658 548 -17624
rect 846 -17658 880 -17624
rect 1012 -17658 1046 -17624
rect 1344 -17658 1378 -17624
rect 1510 -17658 1544 -17624
rect 1842 -17658 1876 -17624
<< psubdiff >>
rect -54 -17792 -30 -17736
rect 1702 -17792 1726 -17736
<< nsubdiff >>
rect -18 -17442 6 -17386
rect 1886 -17442 1910 -17386
<< psubdiffcont >>
rect -30 -17792 1702 -17736
<< nsubdiffcont >>
rect 6 -17442 1886 -17386
<< poly >>
rect -120 -17568 -54 -17552
rect -120 -17602 -104 -17568
rect -70 -17602 -18 -17568
rect 84 -17602 314 -17568
rect 416 -17602 480 -17568
rect 582 -17602 812 -17568
rect 914 -17602 978 -17568
rect 1080 -17602 1310 -17568
rect 1412 -17602 1476 -17568
rect 1578 -17602 1808 -17568
rect 1910 -17602 1936 -17568
rect -120 -17618 -54 -17602
rect -118 -17952 -52 -17936
rect -118 -17986 -102 -17952
rect -68 -17986 978 -17952
rect 1080 -17986 1476 -17952
rect 1578 -17986 1992 -17952
rect -118 -18002 -52 -17986
rect -118 -18094 -52 -18078
rect -118 -18128 -102 -18094
rect -68 -18128 1476 -18094
rect 1578 -18128 1992 -18094
rect -118 -18144 -52 -18128
<< polycont >>
rect -104 -17602 -70 -17568
rect -102 -17986 -68 -17952
rect -102 -18128 -68 -18094
<< locali >>
rect -50 -17386 1942 -17366
rect -50 -17442 6 -17386
rect 1886 -17442 1942 -17386
rect -50 -17462 1942 -17442
rect -18 -17512 84 -17462
rect -18 -17546 -2 -17512
rect 66 -17546 84 -17512
rect -120 -17568 -54 -17552
rect -18 -17562 84 -17546
rect 314 -17512 416 -17462
rect 314 -17546 330 -17512
rect 398 -17546 416 -17512
rect 314 -17562 416 -17546
rect 480 -17512 582 -17462
rect 480 -17546 496 -17512
rect 564 -17546 582 -17512
rect 480 -17562 582 -17546
rect 812 -17512 914 -17462
rect 812 -17546 828 -17512
rect 896 -17546 914 -17512
rect 812 -17562 914 -17546
rect 978 -17512 1080 -17462
rect 978 -17546 994 -17512
rect 1062 -17546 1080 -17512
rect 978 -17562 1080 -17546
rect 1310 -17512 1412 -17462
rect 1310 -17546 1326 -17512
rect 1394 -17546 1412 -17512
rect 1310 -17562 1412 -17546
rect 1476 -17512 1578 -17462
rect 1476 -17546 1492 -17512
rect 1560 -17546 1578 -17512
rect 1476 -17562 1578 -17546
rect 1808 -17512 1910 -17462
rect 1808 -17546 1824 -17512
rect 1892 -17546 1910 -17512
rect 1808 -17562 1910 -17546
rect -120 -17602 -104 -17568
rect -70 -17602 -54 -17568
rect -120 -17716 -54 -17602
rect 0 -17624 66 -17608
rect 0 -17658 16 -17624
rect 50 -17658 66 -17624
rect 0 -17674 66 -17658
rect 332 -17624 398 -17608
rect 332 -17658 348 -17624
rect 382 -17658 398 -17624
rect 332 -17674 398 -17658
rect 498 -17624 564 -17608
rect 498 -17658 514 -17624
rect 548 -17658 564 -17624
rect 498 -17674 564 -17658
rect 830 -17624 896 -17608
rect 830 -17658 846 -17624
rect 880 -17658 896 -17624
rect 830 -17674 896 -17658
rect 996 -17624 1062 -17608
rect 996 -17658 1012 -17624
rect 1046 -17658 1062 -17624
rect 996 -17674 1062 -17658
rect 1328 -17624 1394 -17608
rect 1328 -17658 1344 -17624
rect 1378 -17658 1394 -17624
rect 1328 -17674 1394 -17658
rect 1494 -17624 1560 -17608
rect 1494 -17658 1510 -17624
rect 1544 -17658 1560 -17624
rect 1494 -17674 1560 -17658
rect 1826 -17624 1892 -17608
rect 1826 -17658 1842 -17624
rect 1876 -17658 1892 -17624
rect 1826 -17674 1892 -17658
rect -120 -17736 1726 -17716
rect -120 -17792 -30 -17736
rect 1702 -17792 1726 -17736
rect -120 -17812 1726 -17792
rect 166 -17834 234 -17812
rect 662 -17834 732 -17812
rect 1162 -17834 1230 -17812
rect 0 -17862 66 -17846
rect 0 -17896 16 -17862
rect 50 -17896 66 -17862
rect -118 -17952 -52 -17936
rect -118 -17986 -102 -17952
rect -68 -17986 -52 -17952
rect -118 -18002 -52 -17986
rect -118 -18094 -52 -18078
rect -118 -18128 -102 -18094
rect -68 -18128 -52 -18094
rect -118 -18144 -52 -18128
rect 0 -18236 66 -17896
rect 166 -17883 233 -17834
rect 332 -17862 398 -17846
rect 166 -18236 232 -17883
rect 332 -17896 348 -17862
rect 382 -17896 398 -17862
rect 332 -18236 398 -17896
rect 498 -17862 564 -17846
rect 498 -17896 514 -17862
rect 548 -17896 564 -17862
rect 498 -18236 564 -17896
rect 663 -17909 730 -17834
rect 664 -18236 730 -17909
rect 830 -17862 896 -17846
rect 830 -17896 846 -17862
rect 880 -17896 896 -17862
rect 830 -18236 896 -17896
rect 996 -17862 1062 -17846
rect 996 -17914 1012 -17862
rect 1046 -17914 1062 -17862
rect 996 -18236 1062 -17914
rect 1162 -17885 1229 -17834
rect 1328 -17862 1394 -17846
rect 1162 -18022 1228 -17885
rect 1162 -18056 1178 -18022
rect 1212 -18056 1228 -18022
rect 1162 -18236 1228 -18056
rect 1328 -17896 1344 -17862
rect 1378 -17896 1394 -17862
rect 1328 -18236 1394 -17896
rect 1494 -17862 1560 -17846
rect 1494 -17914 1510 -17862
rect 1544 -17914 1560 -17862
rect 1494 -18164 1560 -17914
rect 1494 -18198 1510 -18164
rect 1544 -18198 1560 -18164
rect 1494 -18236 1560 -18198
rect 1660 -18022 1726 -17812
rect 1660 -18056 1676 -18022
rect 1710 -18056 1726 -18022
rect 1660 -18236 1726 -18056
rect 1826 -17862 1892 -17846
rect 1826 -17896 1842 -17862
rect 1876 -17896 1892 -17862
rect 1826 -18236 1892 -17896
<< viali >>
rect 16 -17658 50 -17624
rect 348 -17658 382 -17624
rect 514 -17658 548 -17624
rect 846 -17658 880 -17624
rect 1012 -17658 1046 -17624
rect 1344 -17658 1378 -17624
rect 1510 -17658 1544 -17624
rect 1842 -17658 1876 -17624
rect 16 -17896 50 -17862
rect 348 -17896 382 -17862
rect 514 -17896 548 -17862
rect 846 -17896 880 -17862
rect 1012 -17880 1046 -17862
rect 1012 -17896 1046 -17880
rect 1344 -17896 1378 -17862
rect 1510 -17880 1544 -17862
rect 1510 -17896 1544 -17880
rect 1842 -17896 1876 -17862
<< metal1 >>
rect 0 -17624 66 -17608
rect 0 -17658 16 -17624
rect 50 -17658 66 -17624
rect 0 -17862 66 -17658
rect 0 -17896 16 -17862
rect 50 -17896 66 -17862
rect 0 -17912 66 -17896
rect 332 -17624 398 -17608
rect 332 -17658 348 -17624
rect 382 -17658 398 -17624
rect 332 -17862 398 -17658
rect 332 -17896 348 -17862
rect 382 -17896 398 -17862
rect 332 -17912 398 -17896
rect 498 -17624 564 -17608
rect 498 -17658 514 -17624
rect 548 -17658 564 -17624
rect 498 -17862 564 -17658
rect 498 -17896 514 -17862
rect 548 -17896 564 -17862
rect 498 -17912 564 -17896
rect 830 -17624 896 -17608
rect 830 -17658 846 -17624
rect 880 -17658 896 -17624
rect 830 -17862 896 -17658
rect 830 -17896 846 -17862
rect 880 -17896 896 -17862
rect 830 -17912 896 -17896
rect 996 -17624 1062 -17608
rect 996 -17658 1012 -17624
rect 1046 -17658 1062 -17624
rect 996 -17862 1062 -17658
rect 996 -17896 1012 -17862
rect 1046 -17896 1062 -17862
rect 996 -17912 1062 -17896
rect 1328 -17624 1394 -17608
rect 1328 -17658 1344 -17624
rect 1378 -17658 1394 -17624
rect 1328 -17862 1394 -17658
rect 1328 -17896 1344 -17862
rect 1378 -17896 1394 -17862
rect 1328 -17912 1394 -17896
rect 1494 -17624 1560 -17608
rect 1494 -17658 1510 -17624
rect 1544 -17658 1560 -17624
rect 1494 -17862 1560 -17658
rect 1494 -17896 1510 -17862
rect 1544 -17896 1560 -17862
rect 1494 -17912 1560 -17896
rect 1826 -17624 1892 -17608
rect 1826 -17658 1842 -17624
rect 1876 -17658 1892 -17624
rect 1826 -17862 1892 -17658
rect 1826 -17896 1842 -17862
rect 1876 -17896 1892 -17862
rect 1826 -17912 1892 -17896
<< labels >>
flabel locali -118 -18002 -52 -17936 0 FreeSerif 160 0 0 0 word126
port 32 nsew
flabel locali -118 -18144 -52 -18078 0 FreeSerif 160 0 0 0 word127
port 35 nsew
flabel locali 332 -18236 398 -18170 0 FreeSerif 160 0 0 0 Y6
port 38 nsew
flabel locali 0 -18236 66 -18170 0 FreeSerif 160 0 0 0 Y7
port 37 nsew
flabel locali 498 -18236 564 -18170 0 FreeSerif 160 0 0 0 Y5
port 39 nsew
flabel locali 830 -18236 896 -18170 0 FreeSerif 160 0 0 0 Y4
port 40 nsew
flabel locali 996 -18236 1062 -18170 0 FreeSerif 160 0 0 0 Y3
port 41 nsew
flabel locali 1328 -18236 1394 -18170 0 FreeSerif 160 0 0 0 Y2
port 42 nsew
flabel locali 1494 -18236 1560 -18170 0 FreeSerif 160 0 0 0 Y1
port 43 nsew
flabel locali 1826 -18236 1892 -18170 0 FreeSerif 160 0 0 0 Y0
port 44 nsew
flabel locali 132 -17812 278 -17716 0 FreeSerif 160 0 0 0 GND!
port 0 nsew
flabel locali -50 -17462 1942 -17366 0 FreeSerif 160 0 0 0 VDD!
port 10 nsew
<< end >>
