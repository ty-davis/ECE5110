magic
tech sky130A
timestamp 1744679307
<< nmos >>
rect -127 -163 -76 -146
rect 5 -234 56 -217
<< ndiff >>
rect -127 -204 56 -171
rect -127 -171 -76 -105
rect 5 -270 56 -204
<< ndiffc >>
rect -110 -130 -93 -113
rect -44 -196 -27 -179
rect 22 -262 39 -245
<< poly >>
rect -381 -163 -127 -146
rect -76 -163 46 -146
rect -381 -234 5 -217
rect 56 -234 69 -217
<< locali >>
rect -118 -113 -85 -105
rect -118 -130 -110 -113
rect -93 -130 -85 -113
rect -118 -270 -85 -130
rect -52 -179 -19 -105
rect -52 -196 -44 -179
rect -27 -196 -19 -179
rect -52 -270 -19 -196
rect 14 -245 47 -105
rect 14 -262 22 -245
rect 39 -262 47 -245
rect 14 -270 47 -262
<< end >>
