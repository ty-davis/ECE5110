magic
tech sky130A
magscale 1 2
timestamp 1745491943
<< error_s >>
rect 60 145672 166 145682
<< nwell >>
rect 7468 150988 7504 151022
<< locali >>
rect 7456 151036 7515 151045
rect 7456 151026 7516 151036
rect 7456 150988 7468 151026
rect 7504 150988 7516 151026
rect 7456 150976 7516 150988
rect 7456 150825 7515 150976
rect 7456 150759 7734 150825
rect 7861 150717 8042 150783
<< viali >>
rect 7468 150988 7504 151026
rect 5687 150757 5757 150827
rect 6083 150783 6137 150837
rect 6317 150765 6371 150819
rect 6719 150783 6773 150837
rect 7067 150685 7121 150739
rect 7175 150685 7229 150739
rect 5268 150623 5322 150677
rect 7414 150658 7480 150724
rect 7807 150717 7861 150783
rect 7580 150558 7622 150594
rect 7888 150554 7928 150596
<< metal1 >>
rect 6435 151103 7632 151169
rect 6435 150907 6501 151103
rect 7450 151035 7521 151041
rect 6549 151026 7521 151035
rect 6549 150988 7468 151026
rect 7504 150988 7521 151026
rect 6549 150976 7521 150988
rect 6070 150843 6150 150850
rect 5674 150833 5770 150840
rect 5674 150751 5681 150833
rect 5763 150751 5770 150833
rect 6070 150777 6077 150843
rect 6143 150777 6150 150843
rect 6070 150770 6150 150777
rect 6304 150825 6384 150832
rect 6304 150759 6311 150825
rect 6377 150759 6384 150825
rect 6304 150752 6384 150759
rect 5674 150744 5770 150751
rect 6549 150709 6608 150976
rect 7450 150970 7521 150976
rect 6707 150777 6713 150843
rect 6779 150777 6785 150843
rect 7061 150739 7127 150751
rect 7061 150685 7067 150739
rect 7121 150685 7127 150739
rect 2268 150607 2352 150618
rect 5256 150617 5262 150683
rect 5328 150617 5334 150683
rect 2251 150604 2352 150607
rect 2251 150552 2268 150604
rect 2342 150552 2352 150604
rect 2251 150541 2317 150552
rect 7061 150409 7127 150685
rect 7169 150739 7235 150751
rect 7169 150685 7175 150739
rect 7229 150685 7235 150739
rect 7169 150513 7235 150685
rect 7402 150730 7492 150738
rect 7402 150652 7408 150730
rect 7486 150652 7492 150730
rect 7402 150644 7492 150652
rect 7566 150594 7632 151103
rect 7801 150783 7867 150795
rect 7566 150558 7580 150594
rect 7622 150558 7632 150594
rect 7566 150542 7632 150558
rect 7759 150717 7807 150783
rect 7861 150717 7867 150783
rect 7759 150705 7867 150717
rect 7759 150513 7825 150705
rect 7169 150447 7825 150513
rect 7874 150596 7940 150608
rect 7874 150554 7888 150596
rect 7928 150554 7940 150596
rect 7874 150409 7940 150554
rect 7061 150343 7940 150409
<< via1 >>
rect 5681 150827 5763 150833
rect 5681 150757 5687 150827
rect 5687 150757 5757 150827
rect 5757 150757 5763 150827
rect 5681 150751 5763 150757
rect 6077 150837 6143 150843
rect 6077 150783 6083 150837
rect 6083 150783 6137 150837
rect 6137 150783 6143 150837
rect 6077 150777 6143 150783
rect 6311 150819 6377 150825
rect 6311 150765 6317 150819
rect 6317 150765 6371 150819
rect 6371 150765 6377 150819
rect 6311 150759 6377 150765
rect 6713 150837 6779 150843
rect 6713 150783 6719 150837
rect 6719 150783 6773 150837
rect 6773 150783 6779 150837
rect 6713 150777 6779 150783
rect 5262 150677 5328 150683
rect 5262 150623 5268 150677
rect 5268 150623 5322 150677
rect 5322 150623 5328 150677
rect 5262 150617 5328 150623
rect -991 150541 -925 150607
rect 2268 150552 2342 150604
rect 7408 150724 7486 150730
rect 7408 150658 7414 150724
rect 7414 150658 7480 150724
rect 7480 150658 7486 150724
rect 7408 150652 7486 150658
<< metal2 >>
rect 6070 150843 6150 150850
rect 5674 150833 5770 150840
rect 5674 150751 5681 150833
rect 5763 150751 5770 150833
rect 6070 150777 6077 150843
rect 6143 150777 6150 150843
rect 6713 150843 6779 150849
rect 6070 150770 6150 150777
rect 6304 150825 6384 150832
rect 6304 150759 6311 150825
rect 6377 150759 6384 150825
rect 6304 150752 6384 150759
rect 5674 150744 5770 150751
rect 5262 150683 5328 150689
rect -1000 150607 -916 150616
rect -6882 150540 -6810 150604
rect -4246 150542 -4148 150606
rect -1000 150541 -991 150607
rect -925 150541 -916 150607
rect 2254 150608 2352 150620
rect 2254 150552 2268 150608
rect 2342 150552 2352 150608
rect 2254 150542 2352 150552
rect 5262 150561 5328 150617
rect 6713 150561 6779 150777
rect 7402 150730 7492 150738
rect 7402 150652 7408 150730
rect 7486 150724 7492 150730
rect 7486 150658 8143 150724
rect 7486 150652 7492 150658
rect 7402 150644 7492 150652
rect -1000 150536 -916 150541
rect 5262 150495 6779 150561
rect 8077 150603 8143 150658
rect 8077 150537 8253 150603
<< via2 >>
rect 5686 150756 5758 150828
rect 6082 150782 6138 150838
rect 6316 150764 6372 150820
rect -991 150541 -925 150607
rect 2268 150604 2342 150608
rect 2268 150552 2342 150604
<< metal3 >>
rect -991 151021 6143 151087
rect -4235 150841 -1273 150923
rect -1193 150841 -1187 150923
rect -4235 150616 -4153 150841
rect -4246 150534 -4148 150616
rect -991 150612 -925 151021
rect -722 150923 -642 150928
rect -723 150922 5763 150923
rect -723 150842 -722 150922
rect -642 150842 5763 150922
rect -723 150841 5763 150842
rect -722 150836 -642 150841
rect 5681 150828 5763 150841
rect 5681 150756 5686 150828
rect 5758 150756 5763 150828
rect 6077 150838 6143 151021
rect 6077 150782 6082 150838
rect 6138 150782 6143 150838
rect 6077 150777 6143 150782
rect 6311 150820 6377 150825
rect 5681 150751 5763 150756
rect 6311 150764 6316 150820
rect 6372 150764 6377 150820
rect 6311 150746 6377 150764
rect -996 150607 -920 150612
rect -996 150541 -991 150607
rect -925 150541 -920 150607
rect 2254 150608 2352 150620
rect 2254 150552 2268 150608
rect 2342 150607 2352 150608
rect 6317 150607 6383 150746
rect 2342 150552 6383 150607
rect 2254 150542 6383 150552
rect 2326 150541 6383 150542
rect -996 150536 -920 150541
<< via3 >>
rect -1273 150841 -1193 150923
rect -722 150842 -642 150922
<< metal4 >>
rect -1274 150923 -1192 150924
rect -1274 150841 -1273 150923
rect -1193 150922 -641 150923
rect -1193 150842 -722 150922
rect -642 150842 -641 150922
rect -1193 150841 -641 150842
rect -1274 150840 -1192 150841
use counter_4  counter_4_0
timestamp 1745485683
transform 1 0 -6640 0 1 150246
box -318 0 12226 976
use counter_8  counter_8_0
timestamp 1745486774
transform 1 0 8428 0 1 150246
box -318 0 25180 976
use decoder_8  decoder_8_0
timestamp 1744679307
transform 1 0 238 0 1 145618
box -238 -145618 5702 1196
use inv  inv_0 ~/magic/library/mag
timestamp 1738780557
transform 1 0 7488 0 1 150246
box -4 0 322 976
use inv  inv_1
timestamp 1738780557
transform 1 0 7796 0 1 150246
box -4 0 322 976
use memory_8  memory_8_0
timestamp 1744679307
transform 1 0 6108 0 1 145480
box -134 -145474 1992 600
use mux4  mux4_0
timestamp 1745483395
transform 1 0 5578 0 1 150246
box 0 0 1914 976
<< labels >>
flabel metal1 7380 151104 7502 151169 0 FreeSerif 160 0 0 0 Freq0
port 2 nsew
flabel metal1 7336 150343 7458 150408 0 FreeSerif 160 0 0 0 Freq1
port 3 nsew
flabel metal2 -6882 150540 -6810 150604 0 FreeSerif 160 0 0 0 CLK
port 1 nsew
<< end >>
