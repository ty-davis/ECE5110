magic
tech sky130A
timestamp 1744679307
<< poly >>
rect 0 -33 33 0
rect 8 -1178 25 -33
rect 66 -33 99 0
rect 74 -1178 91 -33
rect 132 -33 165 0
rect 140 -1178 157 -33
rect 198 -33 231 0
rect 206 -1178 223 -33
rect 264 -33 297 0
rect 272 -1178 289 -33
rect 330 -33 363 0
rect 338 -1178 355 -33
rect 396 -33 429 0
rect 404 -1178 421 -33
rect 462 -33 495 0
rect 470 -1178 487 -33
rect 659 -33 692 0
rect 667 -1178 684 -33
rect 725 -33 758 0
rect 733 -1178 750 -33
rect 791 -33 824 0
rect 799 -1178 816 -33
rect 857 -33 890 0
rect 865 -1178 882 -33
rect 923 -33 956 0
rect 931 -1178 948 -33
rect 989 -33 1022 0
rect 997 -1178 1014 -33
rect 1055 -33 1088 0
rect 1063 -1178 1080 -33
rect 1121 -33 1154 0
rect 1129 -1178 1146 -33
rect 53 142 89 175
rect 36 69 53 248
rect 185 142 221 175
rect 168 69 185 248
rect 317 142 353 175
rect 300 69 317 248
rect 449 142 485 175
rect 432 69 449 248
rect 669 142 705 175
rect 705 69 722 248
rect 801 142 837 175
rect 837 69 854 248
rect 933 142 969 175
rect 969 69 986 248
rect 1065 142 1101 175
rect 1101 69 1118 248
<< polycont >>
rect 8 -25 25 -8
rect 74 -25 91 -8
rect 140 -25 157 -8
rect 206 -25 223 -8
rect 272 -25 289 -8
rect 338 -25 355 -8
rect 404 -25 421 -8
rect 470 -25 487 -8
rect 667 -25 684 -8
rect 733 -25 750 -8
rect 799 -25 816 -8
rect 865 -25 882 -8
rect 931 -25 948 -8
rect 997 -25 1014 -8
rect 1063 -25 1080 -8
rect 1129 -25 1146 -8
rect 64 150 81 167
rect 196 150 213 167
rect 328 150 345 167
rect 460 150 477 167
rect 677 150 694 167
rect 809 150 826 167
rect 941 150 958 167
rect 1073 150 1090 167
<< locali >>
rect 0 -33 33 0
rect 66 -33 99 0
rect 132 -33 165 0
rect 198 -33 231 0
rect 264 -33 297 0
rect 330 -33 363 0
rect 396 -33 429 0
rect 462 -33 495 0
rect 659 -33 692 0
rect 725 -33 758 0
rect 791 -33 824 0
rect 857 -33 890 0
rect 923 -33 956 0
rect 989 -33 1022 0
rect 1055 -33 1088 0
rect 1121 -33 1154 0
rect -53 -100 -33 -57
rect -33 -100 0 -57
rect 33 -100 66 -57
rect 0 -100 33 -57
rect 99 -100 132 -57
rect 165 -100 198 -57
rect 132 -100 165 -57
rect 231 -100 264 -57
rect 297 -100 330 -57
rect 264 -100 297 -57
rect 363 -100 396 -57
rect 429 -100 462 -57
rect 396 -100 429 -57
rect 495 -100 528 -57
rect -53 -171 -33 -128
rect -33 -171 0 -128
rect 33 -171 66 -128
rect 0 -171 33 -128
rect 99 -171 132 -128
rect 165 -171 198 -128
rect 132 -171 165 -128
rect 231 -171 264 -128
rect 297 -171 330 -128
rect 264 -171 297 -128
rect 363 -171 396 -128
rect 429 -171 462 -128
rect 462 -171 495 -128
rect 495 -171 528 -128
rect -53 -242 -33 -199
rect -33 -242 0 -199
rect 33 -242 66 -199
rect 0 -242 33 -199
rect 99 -242 132 -199
rect 165 -242 198 -199
rect 132 -242 165 -199
rect 231 -242 264 -199
rect 297 -242 330 -199
rect 330 -242 363 -199
rect 363 -242 396 -199
rect 429 -242 462 -199
rect 396 -242 429 -199
rect 495 -242 528 -199
rect -53 -313 -33 -270
rect -33 -313 0 -270
rect 33 -313 66 -270
rect 0 -313 33 -270
rect 99 -313 132 -270
rect 165 -313 198 -270
rect 132 -313 165 -270
rect 231 -313 264 -270
rect 297 -313 330 -270
rect 330 -313 363 -270
rect 363 -313 396 -270
rect 429 -313 462 -270
rect 462 -313 495 -270
rect 495 -313 528 -270
rect -53 -384 -33 -341
rect -33 -384 0 -341
rect 33 -384 66 -341
rect 0 -384 33 -341
rect 99 -384 132 -341
rect 165 -384 198 -341
rect 198 -384 231 -341
rect 231 -384 264 -341
rect 297 -384 330 -341
rect 264 -384 297 -341
rect 363 -384 396 -341
rect 429 -384 462 -341
rect 396 -384 429 -341
rect 495 -384 528 -341
rect -53 -455 -33 -412
rect -33 -455 0 -412
rect 33 -455 66 -412
rect 0 -455 33 -412
rect 99 -455 132 -412
rect 165 -455 198 -412
rect 198 -455 231 -412
rect 231 -455 264 -412
rect 297 -455 330 -412
rect 264 -455 297 -412
rect 363 -455 396 -412
rect 429 -455 462 -412
rect 462 -455 495 -412
rect 495 -455 528 -412
rect -53 -526 -33 -483
rect -33 -526 0 -483
rect 33 -526 66 -483
rect 0 -526 33 -483
rect 99 -526 132 -483
rect 165 -526 198 -483
rect 198 -526 231 -483
rect 231 -526 264 -483
rect 297 -526 330 -483
rect 330 -526 363 -483
rect 363 -526 396 -483
rect 429 -526 462 -483
rect 396 -526 429 -483
rect 495 -526 528 -483
rect -53 -597 -33 -554
rect -33 -597 0 -554
rect 33 -597 66 -554
rect 0 -597 33 -554
rect 99 -597 132 -554
rect 165 -597 198 -554
rect 198 -597 231 -554
rect 231 -597 264 -554
rect 297 -597 330 -554
rect 330 -597 363 -554
rect 363 -597 396 -554
rect 429 -597 462 -554
rect 462 -597 495 -554
rect 495 -597 528 -554
rect -53 -668 -33 -625
rect -33 -668 0 -625
rect 33 -668 66 -625
rect 66 -668 99 -625
rect 99 -668 132 -625
rect 165 -668 198 -625
rect 132 -668 165 -625
rect 231 -668 264 -625
rect 297 -668 330 -625
rect 264 -668 297 -625
rect 363 -668 396 -625
rect 429 -668 462 -625
rect 396 -668 429 -625
rect 495 -668 528 -625
rect -53 -739 -33 -696
rect -33 -739 0 -696
rect 33 -739 66 -696
rect 66 -739 99 -696
rect 99 -739 132 -696
rect 165 -739 198 -696
rect 132 -739 165 -696
rect 231 -739 264 -696
rect 297 -739 330 -696
rect 264 -739 297 -696
rect 363 -739 396 -696
rect 429 -739 462 -696
rect 462 -739 495 -696
rect 495 -739 528 -696
rect -53 -810 -33 -767
rect -33 -810 0 -767
rect 33 -810 66 -767
rect 66 -810 99 -767
rect 99 -810 132 -767
rect 165 -810 198 -767
rect 132 -810 165 -767
rect 231 -810 264 -767
rect 297 -810 330 -767
rect 330 -810 363 -767
rect 363 -810 396 -767
rect 429 -810 462 -767
rect 396 -810 429 -767
rect 495 -810 528 -767
rect -53 -881 -33 -838
rect -33 -881 0 -838
rect 33 -881 66 -838
rect 66 -881 99 -838
rect 99 -881 132 -838
rect 165 -881 198 -838
rect 132 -881 165 -838
rect 231 -881 264 -838
rect 297 -881 330 -838
rect 330 -881 363 -838
rect 363 -881 396 -838
rect 429 -881 462 -838
rect 462 -881 495 -838
rect 495 -881 528 -838
rect -53 -952 -33 -909
rect -33 -952 0 -909
rect 33 -952 66 -909
rect 66 -952 99 -909
rect 99 -952 132 -909
rect 165 -952 198 -909
rect 198 -952 231 -909
rect 231 -952 264 -909
rect 297 -952 330 -909
rect 264 -952 297 -909
rect 363 -952 396 -909
rect 429 -952 462 -909
rect 396 -952 429 -909
rect 495 -952 528 -909
rect -53 -1023 -33 -980
rect -33 -1023 0 -980
rect 33 -1023 66 -980
rect 66 -1023 99 -980
rect 99 -1023 132 -980
rect 165 -1023 198 -980
rect 198 -1023 231 -980
rect 231 -1023 264 -980
rect 297 -1023 330 -980
rect 264 -1023 297 -980
rect 363 -1023 396 -980
rect 429 -1023 462 -980
rect 462 -1023 495 -980
rect 495 -1023 528 -980
rect -53 -1094 -33 -1051
rect -33 -1094 0 -1051
rect 33 -1094 66 -1051
rect 66 -1094 99 -1051
rect 99 -1094 132 -1051
rect 165 -1094 198 -1051
rect 198 -1094 231 -1051
rect 231 -1094 264 -1051
rect 297 -1094 330 -1051
rect 330 -1094 363 -1051
rect 363 -1094 396 -1051
rect 429 -1094 462 -1051
rect 396 -1094 429 -1051
rect 495 -1094 528 -1051
rect -53 -1165 -33 -1122
rect -33 -1165 0 -1122
rect 33 -1165 66 -1122
rect 66 -1165 99 -1122
rect 99 -1165 132 -1122
rect 165 -1165 198 -1122
rect 198 -1165 231 -1122
rect 231 -1165 264 -1122
rect 297 -1165 330 -1122
rect 330 -1165 363 -1122
rect 363 -1165 396 -1122
rect 429 -1165 462 -1122
rect 462 -1165 495 -1122
rect 495 -1165 528 -1122
rect 626 -100 659 -57
rect 528 -100 626 -57
rect 626 -100 659 -57
rect 692 -128 725 -57
rect 758 -100 791 -57
rect 824 -128 857 -57
rect 890 -100 923 -57
rect 956 -128 989 -57
rect 1022 -100 1055 -57
rect 1088 -128 1121 -57
rect 626 -171 659 -128
rect 528 -171 626 -128
rect 626 -171 659 -128
rect 692 -199 725 -128
rect 758 -171 791 -128
rect 824 -199 857 -128
rect 890 -171 923 -128
rect 956 -199 989 -128
rect 1022 -171 1055 -128
rect 1088 -199 1121 -128
rect 626 -242 659 -199
rect 528 -242 626 -199
rect 626 -242 659 -199
rect 692 -270 725 -199
rect 758 -242 791 -199
rect 824 -270 857 -199
rect 890 -242 923 -199
rect 956 -270 989 -199
rect 1022 -242 1055 -199
rect 1088 -270 1121 -199
rect 626 -313 659 -270
rect 528 -313 626 -270
rect 626 -313 659 -270
rect 692 -341 725 -270
rect 758 -313 791 -270
rect 824 -341 857 -270
rect 890 -313 923 -270
rect 956 -341 989 -270
rect 1022 -313 1055 -270
rect 1088 -341 1121 -270
rect 626 -384 659 -341
rect 528 -384 626 -341
rect 626 -384 659 -341
rect 692 -412 725 -341
rect 758 -384 791 -341
rect 824 -412 857 -341
rect 890 -384 923 -341
rect 956 -412 989 -341
rect 1022 -384 1055 -341
rect 1088 -412 1121 -341
rect 626 -455 659 -412
rect 528 -455 626 -412
rect 626 -455 659 -412
rect 692 -483 725 -412
rect 758 -455 791 -412
rect 824 -483 857 -412
rect 890 -455 923 -412
rect 956 -483 989 -412
rect 1022 -455 1055 -412
rect 1088 -483 1121 -412
rect 626 -526 659 -483
rect 528 -526 626 -483
rect 626 -526 659 -483
rect 692 -554 725 -483
rect 758 -526 791 -483
rect 824 -554 857 -483
rect 890 -526 923 -483
rect 956 -554 989 -483
rect 1022 -526 1055 -483
rect 1088 -554 1121 -483
rect 626 -597 659 -554
rect 528 -597 626 -554
rect 626 -597 659 -554
rect 692 -625 725 -554
rect 758 -597 791 -554
rect 824 -625 857 -554
rect 890 -597 923 -554
rect 956 -625 989 -554
rect 1022 -597 1055 -554
rect 1088 -625 1121 -554
rect 626 -668 659 -625
rect 528 -668 626 -625
rect 626 -668 659 -625
rect 692 -696 725 -625
rect 758 -668 791 -625
rect 824 -696 857 -625
rect 890 -668 923 -625
rect 956 -696 989 -625
rect 1022 -668 1055 -625
rect 1154 -668 1187 -625
rect 1088 -696 1121 -625
rect 626 -739 659 -696
rect 528 -739 626 -696
rect 626 -739 659 -696
rect 692 -767 725 -696
rect 758 -739 791 -696
rect 824 -767 857 -696
rect 890 -739 923 -696
rect 956 -767 989 -696
rect 1022 -739 1055 -696
rect 1154 -739 1187 -696
rect 1088 -767 1121 -696
rect 626 -810 659 -767
rect 528 -810 626 -767
rect 626 -810 659 -767
rect 692 -838 725 -767
rect 758 -810 791 -767
rect 824 -838 857 -767
rect 890 -810 923 -767
rect 956 -838 989 -767
rect 1022 -810 1055 -767
rect 1154 -810 1187 -767
rect 1088 -838 1121 -767
rect 626 -881 659 -838
rect 528 -881 626 -838
rect 626 -881 659 -838
rect 692 -909 725 -838
rect 758 -881 791 -838
rect 824 -909 857 -838
rect 890 -881 923 -838
rect 956 -909 989 -838
rect 1022 -881 1055 -838
rect 1154 -881 1187 -838
rect 1088 -909 1121 -838
rect 626 -952 659 -909
rect 528 -952 626 -909
rect 626 -952 659 -909
rect 692 -980 725 -909
rect 758 -952 791 -909
rect 824 -980 857 -909
rect 890 -952 923 -909
rect 956 -980 989 -909
rect 1022 -952 1055 -909
rect 1154 -952 1187 -909
rect 1088 -980 1121 -909
rect 626 -1023 659 -980
rect 528 -1023 626 -980
rect 626 -1023 659 -980
rect 692 -1051 725 -980
rect 758 -1023 791 -980
rect 824 -1051 857 -980
rect 890 -1023 923 -980
rect 956 -1051 989 -980
rect 1022 -1023 1055 -980
rect 1154 -1023 1187 -980
rect 1088 -1051 1121 -980
rect 626 -1094 659 -1051
rect 528 -1094 626 -1051
rect 626 -1094 659 -1051
rect 692 -1122 725 -1051
rect 758 -1094 791 -1051
rect 824 -1122 857 -1051
rect 890 -1094 923 -1051
rect 956 -1122 989 -1051
rect 1022 -1094 1055 -1051
rect 1154 -1094 1187 -1051
rect 1088 -1122 1121 -1051
rect 626 -1165 659 -1122
rect 528 -1165 626 -1122
rect 626 -1165 659 -1122
rect 692 -1193 725 -1122
rect 758 -1165 791 -1122
rect 824 -1193 857 -1122
rect 890 -1165 923 -1122
rect 956 -1193 989 -1122
rect 1022 -1165 1055 -1122
rect 1154 -1165 1187 -1122
rect 1088 -1193 1121 -1122
rect -101 17 1154 65
rect -101 252 1154 300
rect -101 -1193 -53 17
rect 626 -1241 1187 -1193
rect 1187 -1241 1267 -1193
rect 1227 -1193 1267 300
rect 1154 252 1227 300
rect 56 65 89 125
rect 0 82 33 125
rect 0 82 33 192
rect 56 142 89 175
rect 0 192 33 235
rect 56 192 89 252
rect 188 65 221 125
rect 132 82 165 125
rect 132 82 165 192
rect 188 142 221 175
rect 132 192 165 235
rect 188 192 221 252
rect 320 65 353 125
rect 264 82 297 125
rect 264 82 297 192
rect 320 142 353 175
rect 264 192 297 235
rect 320 192 353 252
rect 452 65 485 125
rect 396 82 429 125
rect 396 82 429 192
rect 452 142 485 175
rect 396 192 429 235
rect 452 192 485 252
rect 669 65 702 125
rect 725 82 758 125
rect 725 82 758 192
rect 669 142 702 175
rect 725 192 758 235
rect 669 192 702 252
rect 801 65 834 125
rect 857 82 890 125
rect 857 82 890 192
rect 801 142 834 175
rect 857 192 890 235
rect 801 192 834 252
rect 933 65 966 125
rect 989 82 1022 125
rect 989 82 1022 192
rect 933 142 966 175
rect 989 192 1022 235
rect 933 192 966 252
rect 1065 65 1098 125
rect 1121 82 1154 125
rect 1121 82 1154 192
rect 1065 142 1098 175
rect 1121 192 1154 235
rect 1065 192 1098 252
<< nwell >>
rect -119 -1195 546 143
rect 546 7 1156 143
<< viali >>
rect 8 -25 25 -8
rect 74 -25 91 -8
rect 140 -25 157 -8
rect 206 -25 223 -8
rect 272 -25 289 -8
rect 338 -25 355 -8
rect 404 -25 421 -8
rect 470 -25 487 -8
rect 667 -25 684 -8
rect 733 -25 750 -8
rect 799 -25 816 -8
rect 865 -25 882 -8
rect 931 -25 948 -8
rect 997 -25 1014 -8
rect 1063 -25 1080 -8
rect 1129 -25 1146 -8
rect 634 -92 651 -65
rect 634 -92 651 -65
rect 766 -92 783 -65
rect 898 -92 915 -65
rect 1030 -92 1047 -65
rect 634 -163 651 -136
rect 634 -163 651 -136
rect 766 -163 783 -136
rect 898 -163 915 -136
rect 1030 -163 1047 -136
rect 634 -234 651 -207
rect 634 -234 651 -207
rect 766 -234 783 -207
rect 898 -234 915 -207
rect 1030 -234 1047 -207
rect 634 -305 651 -278
rect 634 -305 651 -278
rect 766 -305 783 -278
rect 898 -305 915 -278
rect 1030 -305 1047 -278
rect 634 -376 651 -349
rect 634 -376 651 -349
rect 766 -376 783 -349
rect 898 -376 915 -349
rect 1030 -376 1047 -349
rect 634 -447 651 -420
rect 634 -447 651 -420
rect 766 -447 783 -420
rect 898 -447 915 -420
rect 1030 -447 1047 -420
rect 634 -518 651 -491
rect 634 -518 651 -491
rect 766 -518 783 -491
rect 898 -518 915 -491
rect 1030 -518 1047 -491
rect 634 -589 651 -562
rect 634 -589 651 -562
rect 766 -589 783 -562
rect 898 -589 915 -562
rect 1030 -589 1047 -562
rect 634 -660 651 -633
rect 634 -660 651 -633
rect 766 -660 783 -633
rect 898 -660 915 -633
rect 1030 -660 1047 -633
rect 634 -731 651 -704
rect 634 -731 651 -704
rect 766 -731 783 -704
rect 898 -731 915 -704
rect 1030 -731 1047 -704
rect 634 -802 651 -775
rect 634 -802 651 -775
rect 766 -802 783 -775
rect 898 -802 915 -775
rect 1030 -802 1047 -775
rect 634 -873 651 -846
rect 634 -873 651 -846
rect 766 -873 783 -846
rect 898 -873 915 -846
rect 1030 -873 1047 -846
rect 634 -944 651 -917
rect 634 -944 651 -917
rect 766 -944 783 -917
rect 898 -944 915 -917
rect 1030 -944 1047 -917
rect 634 -1015 651 -988
rect 634 -1015 651 -988
rect 766 -1015 783 -988
rect 898 -1015 915 -988
rect 1030 -1015 1047 -988
rect 634 -1086 651 -1059
rect 634 -1086 651 -1059
rect 766 -1086 783 -1059
rect 898 -1086 915 -1059
rect 1030 -1086 1047 -1059
rect 634 -1157 651 -1130
rect 634 -1157 651 -1130
rect 766 -1157 783 -1130
rect 898 -1157 915 -1130
rect 1030 -1157 1047 -1130
rect 8 90 25 117
rect 64 150 81 167
rect 140 90 157 117
rect 196 150 213 167
rect 272 90 289 117
rect 328 150 345 167
rect 404 90 421 117
rect 460 150 477 167
rect 733 90 750 117
rect 677 150 694 167
rect 865 90 882 117
rect 809 150 826 167
rect 997 90 1014 117
rect 941 150 958 167
rect 1129 90 1146 117
rect 1073 150 1090 167
<< metal1 >>
rect 0 -33 33 0
rect 66 -33 99 0
rect 132 -33 165 0
rect 198 -33 231 0
rect 264 -33 297 0
rect 330 -33 363 0
rect 396 -33 429 0
rect 462 -33 495 0
rect 659 -33 692 0
rect 725 -33 758 0
rect 791 -33 824 0
rect 857 -33 890 0
rect 923 -33 956 0
rect 989 -33 1022 0
rect 1055 -33 1088 0
rect 1121 -33 1154 0
rect 626 -100 1187 -57
rect 626 -171 1187 -128
rect 626 -242 1187 -199
rect 626 -313 1187 -270
rect 626 -384 1187 -341
rect 626 -455 1187 -412
rect 626 -526 1187 -483
rect 626 -597 1187 -554
rect 626 -668 1187 -625
rect 626 -739 1187 -696
rect 626 -810 1187 -767
rect 626 -881 1187 -838
rect 626 -952 1187 -909
rect 626 -1023 1187 -980
rect 626 -1094 1187 -1051
rect 626 -1165 1187 -1122
rect 0 0 33 125
rect 56 142 89 175
rect 66 0 99 175
rect 132 0 165 125
rect 188 142 221 175
rect 198 0 231 175
rect 264 0 297 125
rect 320 142 353 175
rect 330 0 363 175
rect 396 0 429 125
rect 452 142 485 175
rect 462 0 495 175
rect 462 175 495 175
rect 659 175 692 175
rect 495 142 659 175
rect 330 175 363 222
rect 791 175 824 222
rect 363 189 791 222
rect 198 175 231 269
rect 923 175 956 269
rect 231 236 923 269
rect 66 175 99 316
rect 1055 175 1088 316
rect 99 283 1055 316
rect 725 0 758 125
rect 669 142 702 175
rect 659 0 692 175
rect 857 0 890 125
rect 801 142 834 175
rect 791 0 824 175
rect 989 0 1022 125
rect 933 142 966 175
rect 923 0 956 175
rect 1121 0 1154 125
rect 1065 142 1098 175
rect 1055 0 1088 175
<< via1 >>
rect 498 145 525 172
rect 366 192 393 219
rect 234 239 261 266
rect 102 286 129 313
<< metal2 >>
rect 495 142 528 175
rect 363 189 396 222
rect 231 236 264 269
rect 99 283 132 316
<< pdiff >>
rect -33 -100 0 -57
rect 33 -100 66 -57
rect 66 -100 99 -57
rect 99 -100 132 -57
rect 165 -100 198 -57
rect 198 -100 231 -57
rect 231 -100 264 -57
rect 297 -100 330 -57
rect 330 -100 363 -57
rect 363 -100 396 -57
rect 429 -100 462 -57
rect 462 -100 495 -57
rect 495 -100 528 -57
rect -33 -171 0 -128
rect 33 -171 66 -128
rect 66 -171 99 -128
rect 99 -171 132 -128
rect 165 -171 198 -128
rect 198 -171 231 -128
rect 231 -171 264 -128
rect 297 -171 330 -128
rect 330 -171 363 -128
rect 363 -171 396 -128
rect 429 -171 462 -128
rect 396 -171 429 -128
rect 495 -171 528 -128
rect -33 -242 0 -199
rect 33 -242 66 -199
rect 66 -242 99 -199
rect 99 -242 132 -199
rect 165 -242 198 -199
rect 198 -242 231 -199
rect 231 -242 264 -199
rect 297 -242 330 -199
rect 264 -242 297 -199
rect 363 -242 396 -199
rect 429 -242 462 -199
rect 462 -242 495 -199
rect 495 -242 528 -199
rect -33 -313 0 -270
rect 33 -313 66 -270
rect 66 -313 99 -270
rect 99 -313 132 -270
rect 165 -313 198 -270
rect 198 -313 231 -270
rect 231 -313 264 -270
rect 297 -313 330 -270
rect 264 -313 297 -270
rect 363 -313 396 -270
rect 429 -313 462 -270
rect 396 -313 429 -270
rect 495 -313 528 -270
rect -33 -384 0 -341
rect 33 -384 66 -341
rect 66 -384 99 -341
rect 99 -384 132 -341
rect 165 -384 198 -341
rect 132 -384 165 -341
rect 231 -384 264 -341
rect 297 -384 330 -341
rect 330 -384 363 -341
rect 363 -384 396 -341
rect 429 -384 462 -341
rect 462 -384 495 -341
rect 495 -384 528 -341
rect -33 -455 0 -412
rect 33 -455 66 -412
rect 66 -455 99 -412
rect 99 -455 132 -412
rect 165 -455 198 -412
rect 132 -455 165 -412
rect 231 -455 264 -412
rect 297 -455 330 -412
rect 330 -455 363 -412
rect 363 -455 396 -412
rect 429 -455 462 -412
rect 396 -455 429 -412
rect 495 -455 528 -412
rect -33 -526 0 -483
rect 33 -526 66 -483
rect 66 -526 99 -483
rect 99 -526 132 -483
rect 165 -526 198 -483
rect 132 -526 165 -483
rect 231 -526 264 -483
rect 297 -526 330 -483
rect 264 -526 297 -483
rect 363 -526 396 -483
rect 429 -526 462 -483
rect 462 -526 495 -483
rect 495 -526 528 -483
rect -33 -597 0 -554
rect 33 -597 66 -554
rect 66 -597 99 -554
rect 99 -597 132 -554
rect 165 -597 198 -554
rect 132 -597 165 -554
rect 231 -597 264 -554
rect 297 -597 330 -554
rect 264 -597 297 -554
rect 363 -597 396 -554
rect 429 -597 462 -554
rect 396 -597 429 -554
rect 495 -597 528 -554
rect -33 -668 0 -625
rect 33 -668 66 -625
rect 0 -668 33 -625
rect 99 -668 132 -625
rect 165 -668 198 -625
rect 198 -668 231 -625
rect 231 -668 264 -625
rect 297 -668 330 -625
rect 330 -668 363 -625
rect 363 -668 396 -625
rect 429 -668 462 -625
rect 462 -668 495 -625
rect 495 -668 528 -625
rect -33 -739 0 -696
rect 33 -739 66 -696
rect 0 -739 33 -696
rect 99 -739 132 -696
rect 165 -739 198 -696
rect 198 -739 231 -696
rect 231 -739 264 -696
rect 297 -739 330 -696
rect 330 -739 363 -696
rect 363 -739 396 -696
rect 429 -739 462 -696
rect 396 -739 429 -696
rect 495 -739 528 -696
rect -33 -810 0 -767
rect 33 -810 66 -767
rect 0 -810 33 -767
rect 99 -810 132 -767
rect 165 -810 198 -767
rect 198 -810 231 -767
rect 231 -810 264 -767
rect 297 -810 330 -767
rect 264 -810 297 -767
rect 363 -810 396 -767
rect 429 -810 462 -767
rect 462 -810 495 -767
rect 495 -810 528 -767
rect -33 -881 0 -838
rect 33 -881 66 -838
rect 0 -881 33 -838
rect 99 -881 132 -838
rect 165 -881 198 -838
rect 198 -881 231 -838
rect 231 -881 264 -838
rect 297 -881 330 -838
rect 264 -881 297 -838
rect 363 -881 396 -838
rect 429 -881 462 -838
rect 396 -881 429 -838
rect 495 -881 528 -838
rect -33 -952 0 -909
rect 33 -952 66 -909
rect 0 -952 33 -909
rect 99 -952 132 -909
rect 165 -952 198 -909
rect 132 -952 165 -909
rect 231 -952 264 -909
rect 297 -952 330 -909
rect 330 -952 363 -909
rect 363 -952 396 -909
rect 429 -952 462 -909
rect 462 -952 495 -909
rect 495 -952 528 -909
rect -33 -1023 0 -980
rect 33 -1023 66 -980
rect 0 -1023 33 -980
rect 99 -1023 132 -980
rect 165 -1023 198 -980
rect 132 -1023 165 -980
rect 231 -1023 264 -980
rect 297 -1023 330 -980
rect 330 -1023 363 -980
rect 363 -1023 396 -980
rect 429 -1023 462 -980
rect 396 -1023 429 -980
rect 495 -1023 528 -980
rect -33 -1094 0 -1051
rect 33 -1094 66 -1051
rect 0 -1094 33 -1051
rect 99 -1094 132 -1051
rect 165 -1094 198 -1051
rect 132 -1094 165 -1051
rect 231 -1094 264 -1051
rect 297 -1094 330 -1051
rect 264 -1094 297 -1051
rect 363 -1094 396 -1051
rect 429 -1094 462 -1051
rect 462 -1094 495 -1051
rect 495 -1094 528 -1051
rect -33 -1165 0 -1122
rect 33 -1165 66 -1122
rect 0 -1165 33 -1122
rect 99 -1165 132 -1122
rect 165 -1165 198 -1122
rect 132 -1165 165 -1122
rect 231 -1165 264 -1122
rect 297 -1165 330 -1122
rect 264 -1165 297 -1122
rect 363 -1165 396 -1122
rect 429 -1165 462 -1122
rect 396 -1165 429 -1122
rect 495 -1165 528 -1122
rect 56 82 89 125
rect 0 82 56 125
rect 188 82 221 125
rect 132 82 188 125
rect 320 82 353 125
rect 264 82 320 125
rect 452 82 485 125
rect 396 82 452 125
rect 669 82 702 125
rect 702 82 758 125
rect 801 82 834 125
rect 834 82 890 125
rect 933 82 966 125
rect 966 82 1022 125
rect 1065 82 1098 125
rect 1098 82 1154 125
<< ndiff >>
rect 626 -100 659 -57
rect 659 -100 692 -57
rect 692 -100 725 -57
rect 758 -100 791 -57
rect 791 -100 824 -57
rect 824 -100 857 -57
rect 890 -100 923 -57
rect 923 -100 956 -57
rect 956 -100 989 -57
rect 1022 -100 1055 -57
rect 1055 -100 1088 -57
rect 1088 -100 1121 -57
rect 725 -171 758 -128
rect 758 -171 791 -128
rect 692 -171 725 -128
rect 758 -171 791 -128
rect 791 -171 824 -128
rect 824 -171 857 -128
rect 890 -171 923 -128
rect 923 -171 956 -128
rect 956 -171 989 -128
rect 1022 -171 1055 -128
rect 1055 -171 1088 -128
rect 1088 -171 1121 -128
rect 626 -242 659 -199
rect 659 -242 692 -199
rect 692 -242 725 -199
rect 857 -242 890 -199
rect 890 -242 923 -199
rect 824 -242 857 -199
rect 890 -242 923 -199
rect 923 -242 956 -199
rect 956 -242 989 -199
rect 1022 -242 1055 -199
rect 1055 -242 1088 -199
rect 1088 -242 1121 -199
rect 725 -313 758 -270
rect 758 -313 791 -270
rect 692 -313 725 -270
rect 857 -313 890 -270
rect 890 -313 923 -270
rect 824 -313 857 -270
rect 890 -313 923 -270
rect 923 -313 956 -270
rect 956 -313 989 -270
rect 1022 -313 1055 -270
rect 1055 -313 1088 -270
rect 1088 -313 1121 -270
rect 626 -384 659 -341
rect 659 -384 692 -341
rect 692 -384 725 -341
rect 758 -384 791 -341
rect 791 -384 824 -341
rect 824 -384 857 -341
rect 989 -384 1022 -341
rect 1022 -384 1055 -341
rect 956 -384 989 -341
rect 1022 -384 1055 -341
rect 1055 -384 1088 -341
rect 1088 -384 1121 -341
rect 725 -455 758 -412
rect 758 -455 791 -412
rect 692 -455 725 -412
rect 758 -455 791 -412
rect 791 -455 824 -412
rect 824 -455 857 -412
rect 989 -455 1022 -412
rect 1022 -455 1055 -412
rect 956 -455 989 -412
rect 1022 -455 1055 -412
rect 1055 -455 1088 -412
rect 1088 -455 1121 -412
rect 626 -526 659 -483
rect 659 -526 692 -483
rect 692 -526 725 -483
rect 857 -526 890 -483
rect 890 -526 923 -483
rect 824 -526 857 -483
rect 989 -526 1022 -483
rect 1022 -526 1055 -483
rect 956 -526 989 -483
rect 1022 -526 1055 -483
rect 1055 -526 1088 -483
rect 1088 -526 1121 -483
rect 725 -597 758 -554
rect 758 -597 791 -554
rect 692 -597 725 -554
rect 857 -597 890 -554
rect 890 -597 923 -554
rect 824 -597 857 -554
rect 989 -597 1022 -554
rect 1022 -597 1055 -554
rect 956 -597 989 -554
rect 1022 -597 1055 -554
rect 1055 -597 1088 -554
rect 1088 -597 1121 -554
rect 626 -668 659 -625
rect 659 -668 692 -625
rect 692 -668 725 -625
rect 758 -668 791 -625
rect 791 -668 824 -625
rect 824 -668 857 -625
rect 890 -668 923 -625
rect 923 -668 956 -625
rect 956 -668 989 -625
rect 1121 -668 1154 -625
rect 1154 -668 1187 -625
rect 1088 -668 1121 -625
rect 725 -739 758 -696
rect 758 -739 791 -696
rect 692 -739 725 -696
rect 758 -739 791 -696
rect 791 -739 824 -696
rect 824 -739 857 -696
rect 890 -739 923 -696
rect 923 -739 956 -696
rect 956 -739 989 -696
rect 1121 -739 1154 -696
rect 1154 -739 1187 -696
rect 1088 -739 1121 -696
rect 626 -810 659 -767
rect 659 -810 692 -767
rect 692 -810 725 -767
rect 857 -810 890 -767
rect 890 -810 923 -767
rect 824 -810 857 -767
rect 890 -810 923 -767
rect 923 -810 956 -767
rect 956 -810 989 -767
rect 1121 -810 1154 -767
rect 1154 -810 1187 -767
rect 1088 -810 1121 -767
rect 725 -881 758 -838
rect 758 -881 791 -838
rect 692 -881 725 -838
rect 857 -881 890 -838
rect 890 -881 923 -838
rect 824 -881 857 -838
rect 890 -881 923 -838
rect 923 -881 956 -838
rect 956 -881 989 -838
rect 1121 -881 1154 -838
rect 1154 -881 1187 -838
rect 1088 -881 1121 -838
rect 626 -952 659 -909
rect 659 -952 692 -909
rect 692 -952 725 -909
rect 758 -952 791 -909
rect 791 -952 824 -909
rect 824 -952 857 -909
rect 989 -952 1022 -909
rect 1022 -952 1055 -909
rect 956 -952 989 -909
rect 1121 -952 1154 -909
rect 1154 -952 1187 -909
rect 1088 -952 1121 -909
rect 725 -1023 758 -980
rect 758 -1023 791 -980
rect 692 -1023 725 -980
rect 758 -1023 791 -980
rect 791 -1023 824 -980
rect 824 -1023 857 -980
rect 989 -1023 1022 -980
rect 1022 -1023 1055 -980
rect 956 -1023 989 -980
rect 1121 -1023 1154 -980
rect 1154 -1023 1187 -980
rect 1088 -1023 1121 -980
rect 626 -1094 659 -1051
rect 659 -1094 692 -1051
rect 692 -1094 725 -1051
rect 857 -1094 890 -1051
rect 890 -1094 923 -1051
rect 824 -1094 857 -1051
rect 989 -1094 1022 -1051
rect 1022 -1094 1055 -1051
rect 956 -1094 989 -1051
rect 1121 -1094 1154 -1051
rect 1154 -1094 1187 -1051
rect 1088 -1094 1121 -1051
rect 725 -1165 758 -1122
rect 758 -1165 791 -1122
rect 692 -1165 725 -1122
rect 857 -1165 890 -1122
rect 890 -1165 923 -1122
rect 824 -1165 857 -1122
rect 989 -1165 1022 -1122
rect 1022 -1165 1055 -1122
rect 956 -1165 989 -1122
rect 1121 -1165 1154 -1122
rect 1154 -1165 1187 -1122
rect 1088 -1165 1121 -1122
rect 0 192 89 235
rect 132 192 221 235
rect 264 192 353 235
rect 396 192 485 235
rect 669 192 758 235
rect 801 192 890 235
rect 933 192 1022 235
rect 1065 192 1154 235
<< pdiffc >>
rect -25 -92 -8 -65
rect 41 -92 58 -65
rect 107 -92 124 -65
rect 173 -92 190 -65
rect 239 -92 256 -65
rect 305 -92 322 -65
rect 371 -92 388 -65
rect 437 -92 454 -65
rect 503 -92 520 -65
rect -25 -163 -8 -136
rect 41 -163 58 -136
rect 107 -163 124 -136
rect 173 -163 190 -136
rect 239 -163 256 -136
rect 305 -163 322 -136
rect 371 -163 388 -136
rect 437 -163 454 -136
rect 503 -163 520 -136
rect -25 -234 -8 -207
rect 41 -234 58 -207
rect 107 -234 124 -207
rect 173 -234 190 -207
rect 239 -234 256 -207
rect 305 -234 322 -207
rect 371 -234 388 -207
rect 437 -234 454 -207
rect 503 -234 520 -207
rect -25 -305 -8 -278
rect 41 -305 58 -278
rect 107 -305 124 -278
rect 173 -305 190 -278
rect 239 -305 256 -278
rect 305 -305 322 -278
rect 371 -305 388 -278
rect 437 -305 454 -278
rect 503 -305 520 -278
rect -25 -376 -8 -349
rect 41 -376 58 -349
rect 107 -376 124 -349
rect 173 -376 190 -349
rect 239 -376 256 -349
rect 305 -376 322 -349
rect 371 -376 388 -349
rect 437 -376 454 -349
rect 503 -376 520 -349
rect -25 -447 -8 -420
rect 41 -447 58 -420
rect 107 -447 124 -420
rect 173 -447 190 -420
rect 239 -447 256 -420
rect 305 -447 322 -420
rect 371 -447 388 -420
rect 437 -447 454 -420
rect 503 -447 520 -420
rect -25 -518 -8 -491
rect 41 -518 58 -491
rect 107 -518 124 -491
rect 173 -518 190 -491
rect 239 -518 256 -491
rect 305 -518 322 -491
rect 371 -518 388 -491
rect 437 -518 454 -491
rect 503 -518 520 -491
rect -25 -589 -8 -562
rect 41 -589 58 -562
rect 107 -589 124 -562
rect 173 -589 190 -562
rect 239 -589 256 -562
rect 305 -589 322 -562
rect 371 -589 388 -562
rect 437 -589 454 -562
rect 503 -589 520 -562
rect -25 -660 -8 -633
rect 41 -660 58 -633
rect 107 -660 124 -633
rect 173 -660 190 -633
rect 239 -660 256 -633
rect 305 -660 322 -633
rect 371 -660 388 -633
rect 437 -660 454 -633
rect 503 -660 520 -633
rect -25 -731 -8 -704
rect 41 -731 58 -704
rect 107 -731 124 -704
rect 173 -731 190 -704
rect 239 -731 256 -704
rect 305 -731 322 -704
rect 371 -731 388 -704
rect 437 -731 454 -704
rect 503 -731 520 -704
rect -25 -802 -8 -775
rect 41 -802 58 -775
rect 107 -802 124 -775
rect 173 -802 190 -775
rect 239 -802 256 -775
rect 305 -802 322 -775
rect 371 -802 388 -775
rect 437 -802 454 -775
rect 503 -802 520 -775
rect -25 -873 -8 -846
rect 41 -873 58 -846
rect 107 -873 124 -846
rect 173 -873 190 -846
rect 239 -873 256 -846
rect 305 -873 322 -846
rect 371 -873 388 -846
rect 437 -873 454 -846
rect 503 -873 520 -846
rect -25 -944 -8 -917
rect 41 -944 58 -917
rect 107 -944 124 -917
rect 173 -944 190 -917
rect 239 -944 256 -917
rect 305 -944 322 -917
rect 371 -944 388 -917
rect 437 -944 454 -917
rect 503 -944 520 -917
rect -25 -1015 -8 -988
rect 41 -1015 58 -988
rect 107 -1015 124 -988
rect 173 -1015 190 -988
rect 239 -1015 256 -988
rect 305 -1015 322 -988
rect 371 -1015 388 -988
rect 437 -1015 454 -988
rect 503 -1015 520 -988
rect -25 -1086 -8 -1059
rect 41 -1086 58 -1059
rect 107 -1086 124 -1059
rect 173 -1086 190 -1059
rect 239 -1086 256 -1059
rect 305 -1086 322 -1059
rect 371 -1086 388 -1059
rect 437 -1086 454 -1059
rect 503 -1086 520 -1059
rect -25 -1157 -8 -1130
rect 41 -1157 58 -1130
rect 107 -1157 124 -1130
rect 173 -1157 190 -1130
rect 239 -1157 256 -1130
rect 305 -1157 322 -1130
rect 371 -1157 388 -1130
rect 437 -1157 454 -1130
rect 503 -1157 520 -1130
rect 64 90 81 117
rect 8 90 25 117
rect 196 90 213 117
rect 140 90 157 117
rect 328 90 345 117
rect 272 90 289 117
rect 460 90 477 117
rect 404 90 421 117
rect 677 90 694 117
rect 733 90 750 117
rect 809 90 826 117
rect 865 90 882 117
rect 941 90 958 117
rect 997 90 1014 117
rect 1073 90 1090 117
rect 1129 90 1146 117
<< ndiffc >>
rect 634 -92 651 -65
rect 700 -92 717 -65
rect 766 -92 783 -65
rect 832 -92 849 -65
rect 898 -92 915 -65
rect 964 -92 981 -65
rect 1030 -92 1047 -65
rect 1096 -92 1113 -65
rect 700 -163 717 -136
rect 766 -163 783 -136
rect 832 -163 849 -136
rect 898 -163 915 -136
rect 964 -163 981 -136
rect 1030 -163 1047 -136
rect 1096 -163 1113 -136
rect 634 -234 651 -207
rect 700 -234 717 -207
rect 832 -234 849 -207
rect 898 -234 915 -207
rect 964 -234 981 -207
rect 1030 -234 1047 -207
rect 1096 -234 1113 -207
rect 700 -305 717 -278
rect 832 -305 849 -278
rect 898 -305 915 -278
rect 964 -305 981 -278
rect 1030 -305 1047 -278
rect 1096 -305 1113 -278
rect 634 -376 651 -349
rect 700 -376 717 -349
rect 766 -376 783 -349
rect 832 -376 849 -349
rect 964 -376 981 -349
rect 1030 -376 1047 -349
rect 1096 -376 1113 -349
rect 700 -447 717 -420
rect 766 -447 783 -420
rect 832 -447 849 -420
rect 964 -447 981 -420
rect 1030 -447 1047 -420
rect 1096 -447 1113 -420
rect 634 -518 651 -491
rect 700 -518 717 -491
rect 832 -518 849 -491
rect 964 -518 981 -491
rect 1030 -518 1047 -491
rect 1096 -518 1113 -491
rect 700 -589 717 -562
rect 832 -589 849 -562
rect 964 -589 981 -562
rect 1030 -589 1047 -562
rect 1096 -589 1113 -562
rect 634 -660 651 -633
rect 700 -660 717 -633
rect 766 -660 783 -633
rect 832 -660 849 -633
rect 898 -660 915 -633
rect 964 -660 981 -633
rect 1162 -660 1179 -633
rect 1096 -660 1113 -633
rect 700 -731 717 -704
rect 766 -731 783 -704
rect 832 -731 849 -704
rect 898 -731 915 -704
rect 964 -731 981 -704
rect 1162 -731 1179 -704
rect 1096 -731 1113 -704
rect 634 -802 651 -775
rect 700 -802 717 -775
rect 832 -802 849 -775
rect 898 -802 915 -775
rect 964 -802 981 -775
rect 1162 -802 1179 -775
rect 1096 -802 1113 -775
rect 700 -873 717 -846
rect 832 -873 849 -846
rect 898 -873 915 -846
rect 964 -873 981 -846
rect 1162 -873 1179 -846
rect 1096 -873 1113 -846
rect 634 -944 651 -917
rect 700 -944 717 -917
rect 766 -944 783 -917
rect 832 -944 849 -917
rect 964 -944 981 -917
rect 1162 -944 1179 -917
rect 1096 -944 1113 -917
rect 700 -1015 717 -988
rect 766 -1015 783 -988
rect 832 -1015 849 -988
rect 964 -1015 981 -988
rect 1162 -1015 1179 -988
rect 1096 -1015 1113 -988
rect 634 -1086 651 -1059
rect 700 -1086 717 -1059
rect 832 -1086 849 -1059
rect 964 -1086 981 -1059
rect 1162 -1086 1179 -1059
rect 1096 -1086 1113 -1059
rect 700 -1157 717 -1130
rect 832 -1157 849 -1130
rect 964 -1157 981 -1130
rect 1162 -1157 1179 -1130
rect 1096 -1157 1113 -1130
rect 8 200 25 227
rect 64 200 81 227
rect 140 200 157 227
rect 196 200 213 227
rect 272 200 289 227
rect 328 200 345 227
rect 404 200 421 227
rect 460 200 477 227
rect 733 200 750 227
rect 677 200 694 227
rect 865 200 882 227
rect 809 200 826 227
rect 997 200 1014 227
rect 941 200 958 227
rect 1129 200 1146 227
rect 1073 200 1090 227
<< nsubdiff >>
rect -89 27 1142 55
rect -91 -1181 -63 5
<< nsubdiffcont >>
rect -77 27 1130 55
rect -91 -1169 -63 -7
<< psubdiff >>
rect -89 262 1142 290
rect 638 -1231 1175 -1203
<< psubdiffcont >>
rect -77 262 1130 290
rect 650 -1231 1163 -1203
<< labels >>
flabel metal1 1154 -100 1187 -57 0 FreeSerif 160 0 0 0 word0
port 100 nsew
flabel metal1 1154 -171 1187 -128 0 FreeSerif 160 0 0 0 word1
port 101 nsew
flabel metal1 1154 -242 1187 -199 0 FreeSerif 160 0 0 0 word2
port 102 nsew
flabel metal1 1154 -313 1187 -270 0 FreeSerif 160 0 0 0 word3
port 103 nsew
flabel metal1 1154 -384 1187 -341 0 FreeSerif 160 0 0 0 word4
port 104 nsew
flabel metal1 1154 -455 1187 -412 0 FreeSerif 160 0 0 0 word5
port 105 nsew
flabel metal1 1154 -526 1187 -483 0 FreeSerif 160 0 0 0 word6
port 106 nsew
flabel metal1 1154 -597 1187 -554 0 FreeSerif 160 0 0 0 word7
port 107 nsew
flabel metal1 1154 -668 1187 -625 0 FreeSerif 160 0 0 0 word8
port 108 nsew
flabel metal1 1154 -739 1187 -696 0 FreeSerif 160 0 0 0 word9
port 109 nsew
flabel metal1 1154 -810 1187 -767 0 FreeSerif 160 0 0 0 word10
port 110 nsew
flabel metal1 1154 -881 1187 -838 0 FreeSerif 160 0 0 0 word11
port 111 nsew
flabel metal1 1154 -952 1187 -909 0 FreeSerif 160 0 0 0 word12
port 112 nsew
flabel metal1 1154 -1023 1187 -980 0 FreeSerif 160 0 0 0 word13
port 113 nsew
flabel metal1 1154 -1094 1187 -1051 0 FreeSerif 160 0 0 0 word14
port 114 nsew
flabel metal1 1154 -1165 1187 -1122 0 FreeSerif 160 0 0 0 word15
port 115 nsew
flabel locali -101 -1193 -53 17 0 FreeSerif 160 0 0 0 VDD!
port 116 nsew
flabel locali 1227 -1193 1267 300 0 FreeSerif 160 0 0 0 GND!
port 117 nsew
flabel metal2 495 142 528 175 0 FreeSerif 160 0 0 0 A0
port 19 nsew
flabel metal2 363 189 396 222 0 FreeSerif 160 0 0 0 A1
port 20 nsew
flabel metal2 231 236 264 269 0 FreeSerif 160 0 0 0 A2
port 21 nsew
flabel metal2 99 283 132 316 0 FreeSerif 160 0 0 0 A3
port 22 nsew
<< end >>