magic
tech sky130A
timestamp 1739996850
<< nwell >>
rect -2 197 323 488
<< nmos >>
rect 72 113 87 163
rect 126 113 141 163
rect 180 113 195 163
rect 234 113 249 163
<< pmos >>
rect 72 315 87 415
rect 126 315 141 415
rect 180 315 195 415
rect 234 315 249 415
<< ndiff >>
rect 36 113 72 163
rect 87 113 126 163
rect 141 113 180 163
rect 195 113 234 163
rect 249 113 285 163
<< pdiff >>
rect 36 407 72 415
rect 36 323 44 407
rect 61 323 72 407
rect 36 315 72 323
rect 87 407 126 415
rect 87 323 98 407
rect 115 323 126 407
rect 87 315 126 323
rect 141 407 180 415
rect 141 323 152 407
rect 169 323 180 407
rect 141 315 180 323
rect 195 407 234 415
rect 195 323 206 407
rect 223 323 234 407
rect 195 315 234 323
rect 249 407 285 415
rect 249 323 260 407
rect 277 323 285 407
rect 249 315 285 323
<< pdiffc >>
rect 44 323 61 407
rect 98 323 115 407
rect 152 323 169 407
rect 206 323 223 407
rect 260 323 277 407
<< psubdiff >>
rect 0 10 12 38
rect 289 10 301 38
<< nsubdiff >>
rect 16 442 28 470
rect 293 442 305 470
<< psubdiffcont >>
rect 12 10 289 38
<< nsubdiffcont >>
rect 28 442 293 470
<< poly >>
rect 72 415 87 428
rect 126 415 141 428
rect 180 415 195 428
rect 234 415 249 428
rect 72 163 87 315
rect 126 163 141 315
rect 180 163 195 315
rect 234 163 249 315
rect 72 100 87 113
rect 126 100 141 113
rect 180 100 195 113
rect 234 100 249 113
<< locali >>
rect 0 470 321 480
rect 0 442 28 470
rect 293 442 321 470
rect 0 432 321 442
rect 36 407 69 432
rect 36 323 44 407
rect 61 323 69 407
rect 36 315 69 323
rect 90 407 123 415
rect 90 323 98 407
rect 115 323 123 407
rect 90 315 123 323
rect 144 407 177 415
rect 144 323 152 407
rect 169 323 177 407
rect 144 315 177 323
rect 198 407 231 415
rect 198 323 206 407
rect 223 323 231 407
rect 198 315 231 323
rect 252 407 285 432
rect 252 323 260 407
rect 277 323 285 407
rect 252 315 285 323
rect 0 38 301 48
rect 0 10 12 38
rect 289 10 301 38
rect 0 0 301 10
<< labels >>
flabel pdiff 72 365 72 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 141 365 141 365 1 FreeSerif 8 0 0 0 S$
flabel locali 0 432 213 480 0 FreeSerif 80 0 0 0 VDD!
port 2 nsew
flabel locali 0 0 213 48 0 FreeSerif 80 0 0 0 GND!
port 3 nsew
flabel pdiff 195 365 195 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 249 365 249 365 1 FreeSerif 8 0 0 0 S$
<< end >>
