magic
tech sky130A
timestamp 1744679307
<< poly >>
rect 0 -33 33 0
rect 8 -9130 25 -33
rect 66 -33 99 0
rect 74 -9130 91 -33
rect 132 -33 165 0
rect 140 -9130 157 -33
rect 198 -33 231 0
rect 206 -9130 223 -33
rect 264 -33 297 0
rect 272 -9130 289 -33
rect 330 -33 363 0
rect 338 -9130 355 -33
rect 396 -33 429 0
rect 404 -9130 421 -33
rect 462 -33 495 0
rect 470 -9130 487 -33
rect 528 -33 561 0
rect 536 -9130 553 -33
rect 594 -33 627 0
rect 602 -9130 619 -33
rect 660 -33 693 0
rect 668 -9130 685 -33
rect 726 -33 759 0
rect 734 -9130 751 -33
rect 792 -33 825 0
rect 800 -9130 817 -33
rect 858 -33 891 0
rect 866 -9130 883 -33
rect 1055 -33 1088 0
rect 1063 -9130 1080 -33
rect 1121 -33 1154 0
rect 1129 -9130 1146 -33
rect 1187 -33 1220 0
rect 1195 -9130 1212 -33
rect 1253 -33 1286 0
rect 1261 -9130 1278 -33
rect 1319 -33 1352 0
rect 1327 -9130 1344 -33
rect 1385 -33 1418 0
rect 1393 -9130 1410 -33
rect 1451 -33 1484 0
rect 1459 -9130 1476 -33
rect 1517 -33 1550 0
rect 1525 -9130 1542 -33
rect 1583 -33 1616 0
rect 1591 -9130 1608 -33
rect 1649 -33 1682 0
rect 1657 -9130 1674 -33
rect 1715 -33 1748 0
rect 1723 -9130 1740 -33
rect 1781 -33 1814 0
rect 1789 -9130 1806 -33
rect 1847 -33 1880 0
rect 1855 -9130 1872 -33
rect 1913 -33 1946 0
rect 1921 -9130 1938 -33
rect 53 142 89 175
rect 36 69 53 248
rect 185 142 221 175
rect 168 69 185 248
rect 317 142 353 175
rect 300 69 317 248
rect 449 142 485 175
rect 432 69 449 248
rect 581 142 617 175
rect 564 69 581 248
rect 713 142 749 175
rect 696 69 713 248
rect 845 142 881 175
rect 828 69 845 248
rect 1065 142 1101 175
rect 1101 69 1118 248
rect 1197 142 1233 175
rect 1233 69 1250 248
rect 1329 142 1365 175
rect 1365 69 1382 248
rect 1461 142 1497 175
rect 1497 69 1514 248
rect 1593 142 1629 175
rect 1629 69 1646 248
rect 1725 142 1761 175
rect 1761 69 1778 248
rect 1857 142 1893 175
rect 1893 69 1910 248
<< polycont >>
rect 8 -25 25 -8
rect 74 -25 91 -8
rect 140 -25 157 -8
rect 206 -25 223 -8
rect 272 -25 289 -8
rect 338 -25 355 -8
rect 404 -25 421 -8
rect 470 -25 487 -8
rect 536 -25 553 -8
rect 602 -25 619 -8
rect 668 -25 685 -8
rect 734 -25 751 -8
rect 800 -25 817 -8
rect 866 -25 883 -8
rect 1063 -25 1080 -8
rect 1129 -25 1146 -8
rect 1195 -25 1212 -8
rect 1261 -25 1278 -8
rect 1327 -25 1344 -8
rect 1393 -25 1410 -8
rect 1459 -25 1476 -8
rect 1525 -25 1542 -8
rect 1591 -25 1608 -8
rect 1657 -25 1674 -8
rect 1723 -25 1740 -8
rect 1789 -25 1806 -8
rect 1855 -25 1872 -8
rect 1921 -25 1938 -8
rect 64 150 81 167
rect 196 150 213 167
rect 328 150 345 167
rect 460 150 477 167
rect 592 150 609 167
rect 724 150 741 167
rect 856 150 873 167
rect 1073 150 1090 167
rect 1205 150 1222 167
rect 1337 150 1354 167
rect 1469 150 1486 167
rect 1601 150 1618 167
rect 1733 150 1750 167
rect 1865 150 1882 167
<< locali >>
rect 0 -33 33 0
rect 66 -33 99 0
rect 132 -33 165 0
rect 198 -33 231 0
rect 264 -33 297 0
rect 330 -33 363 0
rect 396 -33 429 0
rect 462 -33 495 0
rect 528 -33 561 0
rect 594 -33 627 0
rect 660 -33 693 0
rect 726 -33 759 0
rect 792 -33 825 0
rect 858 -33 891 0
rect 1055 -33 1088 0
rect 1121 -33 1154 0
rect 1187 -33 1220 0
rect 1253 -33 1286 0
rect 1319 -33 1352 0
rect 1385 -33 1418 0
rect 1451 -33 1484 0
rect 1517 -33 1550 0
rect 1583 -33 1616 0
rect 1649 -33 1682 0
rect 1715 -33 1748 0
rect 1781 -33 1814 0
rect 1847 -33 1880 0
rect 1913 -33 1946 0
rect -53 -100 -33 -57
rect -33 -100 0 -57
rect 33 -100 66 -57
rect 0 -100 33 -57
rect 99 -100 132 -57
rect 165 -100 198 -57
rect 132 -100 165 -57
rect 231 -100 264 -57
rect 297 -100 330 -57
rect 264 -100 297 -57
rect 363 -100 396 -57
rect 429 -100 462 -57
rect 396 -100 429 -57
rect 495 -100 528 -57
rect 561 -100 594 -57
rect 528 -100 561 -57
rect 627 -100 660 -57
rect 693 -100 726 -57
rect 660 -100 693 -57
rect 759 -100 792 -57
rect 825 -100 858 -57
rect 792 -100 825 -57
rect 891 -100 924 -57
rect -53 -171 -33 -128
rect -33 -171 0 -128
rect 33 -171 66 -128
rect 0 -171 33 -128
rect 99 -171 132 -128
rect 165 -171 198 -128
rect 132 -171 165 -128
rect 231 -171 264 -128
rect 297 -171 330 -128
rect 264 -171 297 -128
rect 363 -171 396 -128
rect 429 -171 462 -128
rect 396 -171 429 -128
rect 495 -171 528 -128
rect 561 -171 594 -128
rect 528 -171 561 -128
rect 627 -171 660 -128
rect 693 -171 726 -128
rect 660 -171 693 -128
rect 759 -171 792 -128
rect 825 -171 858 -128
rect 858 -171 891 -128
rect 891 -171 924 -128
rect -53 -242 -33 -199
rect -33 -242 0 -199
rect 33 -242 66 -199
rect 0 -242 33 -199
rect 99 -242 132 -199
rect 165 -242 198 -199
rect 132 -242 165 -199
rect 231 -242 264 -199
rect 297 -242 330 -199
rect 264 -242 297 -199
rect 363 -242 396 -199
rect 429 -242 462 -199
rect 396 -242 429 -199
rect 495 -242 528 -199
rect 561 -242 594 -199
rect 528 -242 561 -199
rect 627 -242 660 -199
rect 693 -242 726 -199
rect 726 -242 759 -199
rect 759 -242 792 -199
rect 825 -242 858 -199
rect 792 -242 825 -199
rect 891 -242 924 -199
rect -53 -313 -33 -270
rect -33 -313 0 -270
rect 33 -313 66 -270
rect 0 -313 33 -270
rect 99 -313 132 -270
rect 165 -313 198 -270
rect 132 -313 165 -270
rect 231 -313 264 -270
rect 297 -313 330 -270
rect 264 -313 297 -270
rect 363 -313 396 -270
rect 429 -313 462 -270
rect 396 -313 429 -270
rect 495 -313 528 -270
rect 561 -313 594 -270
rect 528 -313 561 -270
rect 627 -313 660 -270
rect 693 -313 726 -270
rect 726 -313 759 -270
rect 759 -313 792 -270
rect 825 -313 858 -270
rect 858 -313 891 -270
rect 891 -313 924 -270
rect -53 -384 -33 -341
rect -33 -384 0 -341
rect 33 -384 66 -341
rect 0 -384 33 -341
rect 99 -384 132 -341
rect 165 -384 198 -341
rect 132 -384 165 -341
rect 231 -384 264 -341
rect 297 -384 330 -341
rect 264 -384 297 -341
rect 363 -384 396 -341
rect 429 -384 462 -341
rect 396 -384 429 -341
rect 495 -384 528 -341
rect 561 -384 594 -341
rect 594 -384 627 -341
rect 627 -384 660 -341
rect 693 -384 726 -341
rect 660 -384 693 -341
rect 759 -384 792 -341
rect 825 -384 858 -341
rect 792 -384 825 -341
rect 891 -384 924 -341
rect -53 -455 -33 -412
rect -33 -455 0 -412
rect 33 -455 66 -412
rect 0 -455 33 -412
rect 99 -455 132 -412
rect 165 -455 198 -412
rect 132 -455 165 -412
rect 231 -455 264 -412
rect 297 -455 330 -412
rect 264 -455 297 -412
rect 363 -455 396 -412
rect 429 -455 462 -412
rect 396 -455 429 -412
rect 495 -455 528 -412
rect 561 -455 594 -412
rect 594 -455 627 -412
rect 627 -455 660 -412
rect 693 -455 726 -412
rect 660 -455 693 -412
rect 759 -455 792 -412
rect 825 -455 858 -412
rect 858 -455 891 -412
rect 891 -455 924 -412
rect -53 -526 -33 -483
rect -33 -526 0 -483
rect 33 -526 66 -483
rect 0 -526 33 -483
rect 99 -526 132 -483
rect 165 -526 198 -483
rect 132 -526 165 -483
rect 231 -526 264 -483
rect 297 -526 330 -483
rect 264 -526 297 -483
rect 363 -526 396 -483
rect 429 -526 462 -483
rect 396 -526 429 -483
rect 495 -526 528 -483
rect 561 -526 594 -483
rect 594 -526 627 -483
rect 627 -526 660 -483
rect 693 -526 726 -483
rect 726 -526 759 -483
rect 759 -526 792 -483
rect 825 -526 858 -483
rect 792 -526 825 -483
rect 891 -526 924 -483
rect -53 -597 -33 -554
rect -33 -597 0 -554
rect 33 -597 66 -554
rect 0 -597 33 -554
rect 99 -597 132 -554
rect 165 -597 198 -554
rect 132 -597 165 -554
rect 231 -597 264 -554
rect 297 -597 330 -554
rect 264 -597 297 -554
rect 363 -597 396 -554
rect 429 -597 462 -554
rect 396 -597 429 -554
rect 495 -597 528 -554
rect 561 -597 594 -554
rect 594 -597 627 -554
rect 627 -597 660 -554
rect 693 -597 726 -554
rect 726 -597 759 -554
rect 759 -597 792 -554
rect 825 -597 858 -554
rect 858 -597 891 -554
rect 891 -597 924 -554
rect -53 -668 -33 -625
rect -33 -668 0 -625
rect 33 -668 66 -625
rect 0 -668 33 -625
rect 99 -668 132 -625
rect 165 -668 198 -625
rect 132 -668 165 -625
rect 231 -668 264 -625
rect 297 -668 330 -625
rect 264 -668 297 -625
rect 363 -668 396 -625
rect 429 -668 462 -625
rect 462 -668 495 -625
rect 495 -668 528 -625
rect 561 -668 594 -625
rect 528 -668 561 -625
rect 627 -668 660 -625
rect 693 -668 726 -625
rect 660 -668 693 -625
rect 759 -668 792 -625
rect 825 -668 858 -625
rect 792 -668 825 -625
rect 891 -668 924 -625
rect -53 -739 -33 -696
rect -33 -739 0 -696
rect 33 -739 66 -696
rect 0 -739 33 -696
rect 99 -739 132 -696
rect 165 -739 198 -696
rect 132 -739 165 -696
rect 231 -739 264 -696
rect 297 -739 330 -696
rect 264 -739 297 -696
rect 363 -739 396 -696
rect 429 -739 462 -696
rect 462 -739 495 -696
rect 495 -739 528 -696
rect 561 -739 594 -696
rect 528 -739 561 -696
rect 627 -739 660 -696
rect 693 -739 726 -696
rect 660 -739 693 -696
rect 759 -739 792 -696
rect 825 -739 858 -696
rect 858 -739 891 -696
rect 891 -739 924 -696
rect -53 -810 -33 -767
rect -33 -810 0 -767
rect 33 -810 66 -767
rect 0 -810 33 -767
rect 99 -810 132 -767
rect 165 -810 198 -767
rect 132 -810 165 -767
rect 231 -810 264 -767
rect 297 -810 330 -767
rect 264 -810 297 -767
rect 363 -810 396 -767
rect 429 -810 462 -767
rect 462 -810 495 -767
rect 495 -810 528 -767
rect 561 -810 594 -767
rect 528 -810 561 -767
rect 627 -810 660 -767
rect 693 -810 726 -767
rect 726 -810 759 -767
rect 759 -810 792 -767
rect 825 -810 858 -767
rect 792 -810 825 -767
rect 891 -810 924 -767
rect -53 -881 -33 -838
rect -33 -881 0 -838
rect 33 -881 66 -838
rect 0 -881 33 -838
rect 99 -881 132 -838
rect 165 -881 198 -838
rect 132 -881 165 -838
rect 231 -881 264 -838
rect 297 -881 330 -838
rect 264 -881 297 -838
rect 363 -881 396 -838
rect 429 -881 462 -838
rect 462 -881 495 -838
rect 495 -881 528 -838
rect 561 -881 594 -838
rect 528 -881 561 -838
rect 627 -881 660 -838
rect 693 -881 726 -838
rect 726 -881 759 -838
rect 759 -881 792 -838
rect 825 -881 858 -838
rect 858 -881 891 -838
rect 891 -881 924 -838
rect -53 -952 -33 -909
rect -33 -952 0 -909
rect 33 -952 66 -909
rect 0 -952 33 -909
rect 99 -952 132 -909
rect 165 -952 198 -909
rect 132 -952 165 -909
rect 231 -952 264 -909
rect 297 -952 330 -909
rect 264 -952 297 -909
rect 363 -952 396 -909
rect 429 -952 462 -909
rect 462 -952 495 -909
rect 495 -952 528 -909
rect 561 -952 594 -909
rect 594 -952 627 -909
rect 627 -952 660 -909
rect 693 -952 726 -909
rect 660 -952 693 -909
rect 759 -952 792 -909
rect 825 -952 858 -909
rect 792 -952 825 -909
rect 891 -952 924 -909
rect -53 -1023 -33 -980
rect -33 -1023 0 -980
rect 33 -1023 66 -980
rect 0 -1023 33 -980
rect 99 -1023 132 -980
rect 165 -1023 198 -980
rect 132 -1023 165 -980
rect 231 -1023 264 -980
rect 297 -1023 330 -980
rect 264 -1023 297 -980
rect 363 -1023 396 -980
rect 429 -1023 462 -980
rect 462 -1023 495 -980
rect 495 -1023 528 -980
rect 561 -1023 594 -980
rect 594 -1023 627 -980
rect 627 -1023 660 -980
rect 693 -1023 726 -980
rect 660 -1023 693 -980
rect 759 -1023 792 -980
rect 825 -1023 858 -980
rect 858 -1023 891 -980
rect 891 -1023 924 -980
rect -53 -1094 -33 -1051
rect -33 -1094 0 -1051
rect 33 -1094 66 -1051
rect 0 -1094 33 -1051
rect 99 -1094 132 -1051
rect 165 -1094 198 -1051
rect 132 -1094 165 -1051
rect 231 -1094 264 -1051
rect 297 -1094 330 -1051
rect 264 -1094 297 -1051
rect 363 -1094 396 -1051
rect 429 -1094 462 -1051
rect 462 -1094 495 -1051
rect 495 -1094 528 -1051
rect 561 -1094 594 -1051
rect 594 -1094 627 -1051
rect 627 -1094 660 -1051
rect 693 -1094 726 -1051
rect 726 -1094 759 -1051
rect 759 -1094 792 -1051
rect 825 -1094 858 -1051
rect 792 -1094 825 -1051
rect 891 -1094 924 -1051
rect -53 -1165 -33 -1122
rect -33 -1165 0 -1122
rect 33 -1165 66 -1122
rect 0 -1165 33 -1122
rect 99 -1165 132 -1122
rect 165 -1165 198 -1122
rect 132 -1165 165 -1122
rect 231 -1165 264 -1122
rect 297 -1165 330 -1122
rect 264 -1165 297 -1122
rect 363 -1165 396 -1122
rect 429 -1165 462 -1122
rect 462 -1165 495 -1122
rect 495 -1165 528 -1122
rect 561 -1165 594 -1122
rect 594 -1165 627 -1122
rect 627 -1165 660 -1122
rect 693 -1165 726 -1122
rect 726 -1165 759 -1122
rect 759 -1165 792 -1122
rect 825 -1165 858 -1122
rect 858 -1165 891 -1122
rect 891 -1165 924 -1122
rect -53 -1236 -33 -1193
rect -33 -1236 0 -1193
rect 33 -1236 66 -1193
rect 0 -1236 33 -1193
rect 99 -1236 132 -1193
rect 165 -1236 198 -1193
rect 132 -1236 165 -1193
rect 231 -1236 264 -1193
rect 297 -1236 330 -1193
rect 330 -1236 363 -1193
rect 363 -1236 396 -1193
rect 429 -1236 462 -1193
rect 396 -1236 429 -1193
rect 495 -1236 528 -1193
rect 561 -1236 594 -1193
rect 528 -1236 561 -1193
rect 627 -1236 660 -1193
rect 693 -1236 726 -1193
rect 660 -1236 693 -1193
rect 759 -1236 792 -1193
rect 825 -1236 858 -1193
rect 792 -1236 825 -1193
rect 891 -1236 924 -1193
rect -53 -1307 -33 -1264
rect -33 -1307 0 -1264
rect 33 -1307 66 -1264
rect 0 -1307 33 -1264
rect 99 -1307 132 -1264
rect 165 -1307 198 -1264
rect 132 -1307 165 -1264
rect 231 -1307 264 -1264
rect 297 -1307 330 -1264
rect 330 -1307 363 -1264
rect 363 -1307 396 -1264
rect 429 -1307 462 -1264
rect 396 -1307 429 -1264
rect 495 -1307 528 -1264
rect 561 -1307 594 -1264
rect 528 -1307 561 -1264
rect 627 -1307 660 -1264
rect 693 -1307 726 -1264
rect 660 -1307 693 -1264
rect 759 -1307 792 -1264
rect 825 -1307 858 -1264
rect 858 -1307 891 -1264
rect 891 -1307 924 -1264
rect -53 -1378 -33 -1335
rect -33 -1378 0 -1335
rect 33 -1378 66 -1335
rect 0 -1378 33 -1335
rect 99 -1378 132 -1335
rect 165 -1378 198 -1335
rect 132 -1378 165 -1335
rect 231 -1378 264 -1335
rect 297 -1378 330 -1335
rect 330 -1378 363 -1335
rect 363 -1378 396 -1335
rect 429 -1378 462 -1335
rect 396 -1378 429 -1335
rect 495 -1378 528 -1335
rect 561 -1378 594 -1335
rect 528 -1378 561 -1335
rect 627 -1378 660 -1335
rect 693 -1378 726 -1335
rect 726 -1378 759 -1335
rect 759 -1378 792 -1335
rect 825 -1378 858 -1335
rect 792 -1378 825 -1335
rect 891 -1378 924 -1335
rect -53 -1449 -33 -1406
rect -33 -1449 0 -1406
rect 33 -1449 66 -1406
rect 0 -1449 33 -1406
rect 99 -1449 132 -1406
rect 165 -1449 198 -1406
rect 132 -1449 165 -1406
rect 231 -1449 264 -1406
rect 297 -1449 330 -1406
rect 330 -1449 363 -1406
rect 363 -1449 396 -1406
rect 429 -1449 462 -1406
rect 396 -1449 429 -1406
rect 495 -1449 528 -1406
rect 561 -1449 594 -1406
rect 528 -1449 561 -1406
rect 627 -1449 660 -1406
rect 693 -1449 726 -1406
rect 726 -1449 759 -1406
rect 759 -1449 792 -1406
rect 825 -1449 858 -1406
rect 858 -1449 891 -1406
rect 891 -1449 924 -1406
rect -53 -1520 -33 -1477
rect -33 -1520 0 -1477
rect 33 -1520 66 -1477
rect 0 -1520 33 -1477
rect 99 -1520 132 -1477
rect 165 -1520 198 -1477
rect 132 -1520 165 -1477
rect 231 -1520 264 -1477
rect 297 -1520 330 -1477
rect 330 -1520 363 -1477
rect 363 -1520 396 -1477
rect 429 -1520 462 -1477
rect 396 -1520 429 -1477
rect 495 -1520 528 -1477
rect 561 -1520 594 -1477
rect 594 -1520 627 -1477
rect 627 -1520 660 -1477
rect 693 -1520 726 -1477
rect 660 -1520 693 -1477
rect 759 -1520 792 -1477
rect 825 -1520 858 -1477
rect 792 -1520 825 -1477
rect 891 -1520 924 -1477
rect -53 -1591 -33 -1548
rect -33 -1591 0 -1548
rect 33 -1591 66 -1548
rect 0 -1591 33 -1548
rect 99 -1591 132 -1548
rect 165 -1591 198 -1548
rect 132 -1591 165 -1548
rect 231 -1591 264 -1548
rect 297 -1591 330 -1548
rect 330 -1591 363 -1548
rect 363 -1591 396 -1548
rect 429 -1591 462 -1548
rect 396 -1591 429 -1548
rect 495 -1591 528 -1548
rect 561 -1591 594 -1548
rect 594 -1591 627 -1548
rect 627 -1591 660 -1548
rect 693 -1591 726 -1548
rect 660 -1591 693 -1548
rect 759 -1591 792 -1548
rect 825 -1591 858 -1548
rect 858 -1591 891 -1548
rect 891 -1591 924 -1548
rect -53 -1662 -33 -1619
rect -33 -1662 0 -1619
rect 33 -1662 66 -1619
rect 0 -1662 33 -1619
rect 99 -1662 132 -1619
rect 165 -1662 198 -1619
rect 132 -1662 165 -1619
rect 231 -1662 264 -1619
rect 297 -1662 330 -1619
rect 330 -1662 363 -1619
rect 363 -1662 396 -1619
rect 429 -1662 462 -1619
rect 396 -1662 429 -1619
rect 495 -1662 528 -1619
rect 561 -1662 594 -1619
rect 594 -1662 627 -1619
rect 627 -1662 660 -1619
rect 693 -1662 726 -1619
rect 726 -1662 759 -1619
rect 759 -1662 792 -1619
rect 825 -1662 858 -1619
rect 792 -1662 825 -1619
rect 891 -1662 924 -1619
rect -53 -1733 -33 -1690
rect -33 -1733 0 -1690
rect 33 -1733 66 -1690
rect 0 -1733 33 -1690
rect 99 -1733 132 -1690
rect 165 -1733 198 -1690
rect 132 -1733 165 -1690
rect 231 -1733 264 -1690
rect 297 -1733 330 -1690
rect 330 -1733 363 -1690
rect 363 -1733 396 -1690
rect 429 -1733 462 -1690
rect 396 -1733 429 -1690
rect 495 -1733 528 -1690
rect 561 -1733 594 -1690
rect 594 -1733 627 -1690
rect 627 -1733 660 -1690
rect 693 -1733 726 -1690
rect 726 -1733 759 -1690
rect 759 -1733 792 -1690
rect 825 -1733 858 -1690
rect 858 -1733 891 -1690
rect 891 -1733 924 -1690
rect -53 -1804 -33 -1761
rect -33 -1804 0 -1761
rect 33 -1804 66 -1761
rect 0 -1804 33 -1761
rect 99 -1804 132 -1761
rect 165 -1804 198 -1761
rect 132 -1804 165 -1761
rect 231 -1804 264 -1761
rect 297 -1804 330 -1761
rect 330 -1804 363 -1761
rect 363 -1804 396 -1761
rect 429 -1804 462 -1761
rect 462 -1804 495 -1761
rect 495 -1804 528 -1761
rect 561 -1804 594 -1761
rect 528 -1804 561 -1761
rect 627 -1804 660 -1761
rect 693 -1804 726 -1761
rect 660 -1804 693 -1761
rect 759 -1804 792 -1761
rect 825 -1804 858 -1761
rect 792 -1804 825 -1761
rect 891 -1804 924 -1761
rect -53 -1875 -33 -1832
rect -33 -1875 0 -1832
rect 33 -1875 66 -1832
rect 0 -1875 33 -1832
rect 99 -1875 132 -1832
rect 165 -1875 198 -1832
rect 132 -1875 165 -1832
rect 231 -1875 264 -1832
rect 297 -1875 330 -1832
rect 330 -1875 363 -1832
rect 363 -1875 396 -1832
rect 429 -1875 462 -1832
rect 462 -1875 495 -1832
rect 495 -1875 528 -1832
rect 561 -1875 594 -1832
rect 528 -1875 561 -1832
rect 627 -1875 660 -1832
rect 693 -1875 726 -1832
rect 660 -1875 693 -1832
rect 759 -1875 792 -1832
rect 825 -1875 858 -1832
rect 858 -1875 891 -1832
rect 891 -1875 924 -1832
rect -53 -1946 -33 -1903
rect -33 -1946 0 -1903
rect 33 -1946 66 -1903
rect 0 -1946 33 -1903
rect 99 -1946 132 -1903
rect 165 -1946 198 -1903
rect 132 -1946 165 -1903
rect 231 -1946 264 -1903
rect 297 -1946 330 -1903
rect 330 -1946 363 -1903
rect 363 -1946 396 -1903
rect 429 -1946 462 -1903
rect 462 -1946 495 -1903
rect 495 -1946 528 -1903
rect 561 -1946 594 -1903
rect 528 -1946 561 -1903
rect 627 -1946 660 -1903
rect 693 -1946 726 -1903
rect 726 -1946 759 -1903
rect 759 -1946 792 -1903
rect 825 -1946 858 -1903
rect 792 -1946 825 -1903
rect 891 -1946 924 -1903
rect -53 -2017 -33 -1974
rect -33 -2017 0 -1974
rect 33 -2017 66 -1974
rect 0 -2017 33 -1974
rect 99 -2017 132 -1974
rect 165 -2017 198 -1974
rect 132 -2017 165 -1974
rect 231 -2017 264 -1974
rect 297 -2017 330 -1974
rect 330 -2017 363 -1974
rect 363 -2017 396 -1974
rect 429 -2017 462 -1974
rect 462 -2017 495 -1974
rect 495 -2017 528 -1974
rect 561 -2017 594 -1974
rect 528 -2017 561 -1974
rect 627 -2017 660 -1974
rect 693 -2017 726 -1974
rect 726 -2017 759 -1974
rect 759 -2017 792 -1974
rect 825 -2017 858 -1974
rect 858 -2017 891 -1974
rect 891 -2017 924 -1974
rect -53 -2088 -33 -2045
rect -33 -2088 0 -2045
rect 33 -2088 66 -2045
rect 0 -2088 33 -2045
rect 99 -2088 132 -2045
rect 165 -2088 198 -2045
rect 132 -2088 165 -2045
rect 231 -2088 264 -2045
rect 297 -2088 330 -2045
rect 330 -2088 363 -2045
rect 363 -2088 396 -2045
rect 429 -2088 462 -2045
rect 462 -2088 495 -2045
rect 495 -2088 528 -2045
rect 561 -2088 594 -2045
rect 594 -2088 627 -2045
rect 627 -2088 660 -2045
rect 693 -2088 726 -2045
rect 660 -2088 693 -2045
rect 759 -2088 792 -2045
rect 825 -2088 858 -2045
rect 792 -2088 825 -2045
rect 891 -2088 924 -2045
rect -53 -2159 -33 -2116
rect -33 -2159 0 -2116
rect 33 -2159 66 -2116
rect 0 -2159 33 -2116
rect 99 -2159 132 -2116
rect 165 -2159 198 -2116
rect 132 -2159 165 -2116
rect 231 -2159 264 -2116
rect 297 -2159 330 -2116
rect 330 -2159 363 -2116
rect 363 -2159 396 -2116
rect 429 -2159 462 -2116
rect 462 -2159 495 -2116
rect 495 -2159 528 -2116
rect 561 -2159 594 -2116
rect 594 -2159 627 -2116
rect 627 -2159 660 -2116
rect 693 -2159 726 -2116
rect 660 -2159 693 -2116
rect 759 -2159 792 -2116
rect 825 -2159 858 -2116
rect 858 -2159 891 -2116
rect 891 -2159 924 -2116
rect -53 -2230 -33 -2187
rect -33 -2230 0 -2187
rect 33 -2230 66 -2187
rect 0 -2230 33 -2187
rect 99 -2230 132 -2187
rect 165 -2230 198 -2187
rect 132 -2230 165 -2187
rect 231 -2230 264 -2187
rect 297 -2230 330 -2187
rect 330 -2230 363 -2187
rect 363 -2230 396 -2187
rect 429 -2230 462 -2187
rect 462 -2230 495 -2187
rect 495 -2230 528 -2187
rect 561 -2230 594 -2187
rect 594 -2230 627 -2187
rect 627 -2230 660 -2187
rect 693 -2230 726 -2187
rect 726 -2230 759 -2187
rect 759 -2230 792 -2187
rect 825 -2230 858 -2187
rect 792 -2230 825 -2187
rect 891 -2230 924 -2187
rect -53 -2301 -33 -2258
rect -33 -2301 0 -2258
rect 33 -2301 66 -2258
rect 0 -2301 33 -2258
rect 99 -2301 132 -2258
rect 165 -2301 198 -2258
rect 132 -2301 165 -2258
rect 231 -2301 264 -2258
rect 297 -2301 330 -2258
rect 330 -2301 363 -2258
rect 363 -2301 396 -2258
rect 429 -2301 462 -2258
rect 462 -2301 495 -2258
rect 495 -2301 528 -2258
rect 561 -2301 594 -2258
rect 594 -2301 627 -2258
rect 627 -2301 660 -2258
rect 693 -2301 726 -2258
rect 726 -2301 759 -2258
rect 759 -2301 792 -2258
rect 825 -2301 858 -2258
rect 858 -2301 891 -2258
rect 891 -2301 924 -2258
rect -53 -2372 -33 -2329
rect -33 -2372 0 -2329
rect 33 -2372 66 -2329
rect 0 -2372 33 -2329
rect 99 -2372 132 -2329
rect 165 -2372 198 -2329
rect 198 -2372 231 -2329
rect 231 -2372 264 -2329
rect 297 -2372 330 -2329
rect 264 -2372 297 -2329
rect 363 -2372 396 -2329
rect 429 -2372 462 -2329
rect 396 -2372 429 -2329
rect 495 -2372 528 -2329
rect 561 -2372 594 -2329
rect 528 -2372 561 -2329
rect 627 -2372 660 -2329
rect 693 -2372 726 -2329
rect 660 -2372 693 -2329
rect 759 -2372 792 -2329
rect 825 -2372 858 -2329
rect 792 -2372 825 -2329
rect 891 -2372 924 -2329
rect -53 -2443 -33 -2400
rect -33 -2443 0 -2400
rect 33 -2443 66 -2400
rect 0 -2443 33 -2400
rect 99 -2443 132 -2400
rect 165 -2443 198 -2400
rect 198 -2443 231 -2400
rect 231 -2443 264 -2400
rect 297 -2443 330 -2400
rect 264 -2443 297 -2400
rect 363 -2443 396 -2400
rect 429 -2443 462 -2400
rect 396 -2443 429 -2400
rect 495 -2443 528 -2400
rect 561 -2443 594 -2400
rect 528 -2443 561 -2400
rect 627 -2443 660 -2400
rect 693 -2443 726 -2400
rect 660 -2443 693 -2400
rect 759 -2443 792 -2400
rect 825 -2443 858 -2400
rect 858 -2443 891 -2400
rect 891 -2443 924 -2400
rect -53 -2514 -33 -2471
rect -33 -2514 0 -2471
rect 33 -2514 66 -2471
rect 0 -2514 33 -2471
rect 99 -2514 132 -2471
rect 165 -2514 198 -2471
rect 198 -2514 231 -2471
rect 231 -2514 264 -2471
rect 297 -2514 330 -2471
rect 264 -2514 297 -2471
rect 363 -2514 396 -2471
rect 429 -2514 462 -2471
rect 396 -2514 429 -2471
rect 495 -2514 528 -2471
rect 561 -2514 594 -2471
rect 528 -2514 561 -2471
rect 627 -2514 660 -2471
rect 693 -2514 726 -2471
rect 726 -2514 759 -2471
rect 759 -2514 792 -2471
rect 825 -2514 858 -2471
rect 792 -2514 825 -2471
rect 891 -2514 924 -2471
rect -53 -2585 -33 -2542
rect -33 -2585 0 -2542
rect 33 -2585 66 -2542
rect 0 -2585 33 -2542
rect 99 -2585 132 -2542
rect 165 -2585 198 -2542
rect 198 -2585 231 -2542
rect 231 -2585 264 -2542
rect 297 -2585 330 -2542
rect 264 -2585 297 -2542
rect 363 -2585 396 -2542
rect 429 -2585 462 -2542
rect 396 -2585 429 -2542
rect 495 -2585 528 -2542
rect 561 -2585 594 -2542
rect 528 -2585 561 -2542
rect 627 -2585 660 -2542
rect 693 -2585 726 -2542
rect 726 -2585 759 -2542
rect 759 -2585 792 -2542
rect 825 -2585 858 -2542
rect 858 -2585 891 -2542
rect 891 -2585 924 -2542
rect -53 -2656 -33 -2613
rect -33 -2656 0 -2613
rect 33 -2656 66 -2613
rect 0 -2656 33 -2613
rect 99 -2656 132 -2613
rect 165 -2656 198 -2613
rect 198 -2656 231 -2613
rect 231 -2656 264 -2613
rect 297 -2656 330 -2613
rect 264 -2656 297 -2613
rect 363 -2656 396 -2613
rect 429 -2656 462 -2613
rect 396 -2656 429 -2613
rect 495 -2656 528 -2613
rect 561 -2656 594 -2613
rect 594 -2656 627 -2613
rect 627 -2656 660 -2613
rect 693 -2656 726 -2613
rect 660 -2656 693 -2613
rect 759 -2656 792 -2613
rect 825 -2656 858 -2613
rect 792 -2656 825 -2613
rect 891 -2656 924 -2613
rect -53 -2727 -33 -2684
rect -33 -2727 0 -2684
rect 33 -2727 66 -2684
rect 0 -2727 33 -2684
rect 99 -2727 132 -2684
rect 165 -2727 198 -2684
rect 198 -2727 231 -2684
rect 231 -2727 264 -2684
rect 297 -2727 330 -2684
rect 264 -2727 297 -2684
rect 363 -2727 396 -2684
rect 429 -2727 462 -2684
rect 396 -2727 429 -2684
rect 495 -2727 528 -2684
rect 561 -2727 594 -2684
rect 594 -2727 627 -2684
rect 627 -2727 660 -2684
rect 693 -2727 726 -2684
rect 660 -2727 693 -2684
rect 759 -2727 792 -2684
rect 825 -2727 858 -2684
rect 858 -2727 891 -2684
rect 891 -2727 924 -2684
rect -53 -2798 -33 -2755
rect -33 -2798 0 -2755
rect 33 -2798 66 -2755
rect 0 -2798 33 -2755
rect 99 -2798 132 -2755
rect 165 -2798 198 -2755
rect 198 -2798 231 -2755
rect 231 -2798 264 -2755
rect 297 -2798 330 -2755
rect 264 -2798 297 -2755
rect 363 -2798 396 -2755
rect 429 -2798 462 -2755
rect 396 -2798 429 -2755
rect 495 -2798 528 -2755
rect 561 -2798 594 -2755
rect 594 -2798 627 -2755
rect 627 -2798 660 -2755
rect 693 -2798 726 -2755
rect 726 -2798 759 -2755
rect 759 -2798 792 -2755
rect 825 -2798 858 -2755
rect 792 -2798 825 -2755
rect 891 -2798 924 -2755
rect -53 -2869 -33 -2826
rect -33 -2869 0 -2826
rect 33 -2869 66 -2826
rect 0 -2869 33 -2826
rect 99 -2869 132 -2826
rect 165 -2869 198 -2826
rect 198 -2869 231 -2826
rect 231 -2869 264 -2826
rect 297 -2869 330 -2826
rect 264 -2869 297 -2826
rect 363 -2869 396 -2826
rect 429 -2869 462 -2826
rect 396 -2869 429 -2826
rect 495 -2869 528 -2826
rect 561 -2869 594 -2826
rect 594 -2869 627 -2826
rect 627 -2869 660 -2826
rect 693 -2869 726 -2826
rect 726 -2869 759 -2826
rect 759 -2869 792 -2826
rect 825 -2869 858 -2826
rect 858 -2869 891 -2826
rect 891 -2869 924 -2826
rect -53 -2940 -33 -2897
rect -33 -2940 0 -2897
rect 33 -2940 66 -2897
rect 0 -2940 33 -2897
rect 99 -2940 132 -2897
rect 165 -2940 198 -2897
rect 198 -2940 231 -2897
rect 231 -2940 264 -2897
rect 297 -2940 330 -2897
rect 264 -2940 297 -2897
rect 363 -2940 396 -2897
rect 429 -2940 462 -2897
rect 462 -2940 495 -2897
rect 495 -2940 528 -2897
rect 561 -2940 594 -2897
rect 528 -2940 561 -2897
rect 627 -2940 660 -2897
rect 693 -2940 726 -2897
rect 660 -2940 693 -2897
rect 759 -2940 792 -2897
rect 825 -2940 858 -2897
rect 792 -2940 825 -2897
rect 891 -2940 924 -2897
rect -53 -3011 -33 -2968
rect -33 -3011 0 -2968
rect 33 -3011 66 -2968
rect 0 -3011 33 -2968
rect 99 -3011 132 -2968
rect 165 -3011 198 -2968
rect 198 -3011 231 -2968
rect 231 -3011 264 -2968
rect 297 -3011 330 -2968
rect 264 -3011 297 -2968
rect 363 -3011 396 -2968
rect 429 -3011 462 -2968
rect 462 -3011 495 -2968
rect 495 -3011 528 -2968
rect 561 -3011 594 -2968
rect 528 -3011 561 -2968
rect 627 -3011 660 -2968
rect 693 -3011 726 -2968
rect 660 -3011 693 -2968
rect 759 -3011 792 -2968
rect 825 -3011 858 -2968
rect 858 -3011 891 -2968
rect 891 -3011 924 -2968
rect -53 -3082 -33 -3039
rect -33 -3082 0 -3039
rect 33 -3082 66 -3039
rect 0 -3082 33 -3039
rect 99 -3082 132 -3039
rect 165 -3082 198 -3039
rect 198 -3082 231 -3039
rect 231 -3082 264 -3039
rect 297 -3082 330 -3039
rect 264 -3082 297 -3039
rect 363 -3082 396 -3039
rect 429 -3082 462 -3039
rect 462 -3082 495 -3039
rect 495 -3082 528 -3039
rect 561 -3082 594 -3039
rect 528 -3082 561 -3039
rect 627 -3082 660 -3039
rect 693 -3082 726 -3039
rect 726 -3082 759 -3039
rect 759 -3082 792 -3039
rect 825 -3082 858 -3039
rect 792 -3082 825 -3039
rect 891 -3082 924 -3039
rect -53 -3153 -33 -3110
rect -33 -3153 0 -3110
rect 33 -3153 66 -3110
rect 0 -3153 33 -3110
rect 99 -3153 132 -3110
rect 165 -3153 198 -3110
rect 198 -3153 231 -3110
rect 231 -3153 264 -3110
rect 297 -3153 330 -3110
rect 264 -3153 297 -3110
rect 363 -3153 396 -3110
rect 429 -3153 462 -3110
rect 462 -3153 495 -3110
rect 495 -3153 528 -3110
rect 561 -3153 594 -3110
rect 528 -3153 561 -3110
rect 627 -3153 660 -3110
rect 693 -3153 726 -3110
rect 726 -3153 759 -3110
rect 759 -3153 792 -3110
rect 825 -3153 858 -3110
rect 858 -3153 891 -3110
rect 891 -3153 924 -3110
rect -53 -3224 -33 -3181
rect -33 -3224 0 -3181
rect 33 -3224 66 -3181
rect 0 -3224 33 -3181
rect 99 -3224 132 -3181
rect 165 -3224 198 -3181
rect 198 -3224 231 -3181
rect 231 -3224 264 -3181
rect 297 -3224 330 -3181
rect 264 -3224 297 -3181
rect 363 -3224 396 -3181
rect 429 -3224 462 -3181
rect 462 -3224 495 -3181
rect 495 -3224 528 -3181
rect 561 -3224 594 -3181
rect 594 -3224 627 -3181
rect 627 -3224 660 -3181
rect 693 -3224 726 -3181
rect 660 -3224 693 -3181
rect 759 -3224 792 -3181
rect 825 -3224 858 -3181
rect 792 -3224 825 -3181
rect 891 -3224 924 -3181
rect -53 -3295 -33 -3252
rect -33 -3295 0 -3252
rect 33 -3295 66 -3252
rect 0 -3295 33 -3252
rect 99 -3295 132 -3252
rect 165 -3295 198 -3252
rect 198 -3295 231 -3252
rect 231 -3295 264 -3252
rect 297 -3295 330 -3252
rect 264 -3295 297 -3252
rect 363 -3295 396 -3252
rect 429 -3295 462 -3252
rect 462 -3295 495 -3252
rect 495 -3295 528 -3252
rect 561 -3295 594 -3252
rect 594 -3295 627 -3252
rect 627 -3295 660 -3252
rect 693 -3295 726 -3252
rect 660 -3295 693 -3252
rect 759 -3295 792 -3252
rect 825 -3295 858 -3252
rect 858 -3295 891 -3252
rect 891 -3295 924 -3252
rect -53 -3366 -33 -3323
rect -33 -3366 0 -3323
rect 33 -3366 66 -3323
rect 0 -3366 33 -3323
rect 99 -3366 132 -3323
rect 165 -3366 198 -3323
rect 198 -3366 231 -3323
rect 231 -3366 264 -3323
rect 297 -3366 330 -3323
rect 264 -3366 297 -3323
rect 363 -3366 396 -3323
rect 429 -3366 462 -3323
rect 462 -3366 495 -3323
rect 495 -3366 528 -3323
rect 561 -3366 594 -3323
rect 594 -3366 627 -3323
rect 627 -3366 660 -3323
rect 693 -3366 726 -3323
rect 726 -3366 759 -3323
rect 759 -3366 792 -3323
rect 825 -3366 858 -3323
rect 792 -3366 825 -3323
rect 891 -3366 924 -3323
rect -53 -3437 -33 -3394
rect -33 -3437 0 -3394
rect 33 -3437 66 -3394
rect 0 -3437 33 -3394
rect 99 -3437 132 -3394
rect 165 -3437 198 -3394
rect 198 -3437 231 -3394
rect 231 -3437 264 -3394
rect 297 -3437 330 -3394
rect 264 -3437 297 -3394
rect 363 -3437 396 -3394
rect 429 -3437 462 -3394
rect 462 -3437 495 -3394
rect 495 -3437 528 -3394
rect 561 -3437 594 -3394
rect 594 -3437 627 -3394
rect 627 -3437 660 -3394
rect 693 -3437 726 -3394
rect 726 -3437 759 -3394
rect 759 -3437 792 -3394
rect 825 -3437 858 -3394
rect 858 -3437 891 -3394
rect 891 -3437 924 -3394
rect -53 -3508 -33 -3465
rect -33 -3508 0 -3465
rect 33 -3508 66 -3465
rect 0 -3508 33 -3465
rect 99 -3508 132 -3465
rect 165 -3508 198 -3465
rect 198 -3508 231 -3465
rect 231 -3508 264 -3465
rect 297 -3508 330 -3465
rect 330 -3508 363 -3465
rect 363 -3508 396 -3465
rect 429 -3508 462 -3465
rect 396 -3508 429 -3465
rect 495 -3508 528 -3465
rect 561 -3508 594 -3465
rect 528 -3508 561 -3465
rect 627 -3508 660 -3465
rect 693 -3508 726 -3465
rect 660 -3508 693 -3465
rect 759 -3508 792 -3465
rect 825 -3508 858 -3465
rect 792 -3508 825 -3465
rect 891 -3508 924 -3465
rect -53 -3579 -33 -3536
rect -33 -3579 0 -3536
rect 33 -3579 66 -3536
rect 0 -3579 33 -3536
rect 99 -3579 132 -3536
rect 165 -3579 198 -3536
rect 198 -3579 231 -3536
rect 231 -3579 264 -3536
rect 297 -3579 330 -3536
rect 330 -3579 363 -3536
rect 363 -3579 396 -3536
rect 429 -3579 462 -3536
rect 396 -3579 429 -3536
rect 495 -3579 528 -3536
rect 561 -3579 594 -3536
rect 528 -3579 561 -3536
rect 627 -3579 660 -3536
rect 693 -3579 726 -3536
rect 660 -3579 693 -3536
rect 759 -3579 792 -3536
rect 825 -3579 858 -3536
rect 858 -3579 891 -3536
rect 891 -3579 924 -3536
rect -53 -3650 -33 -3607
rect -33 -3650 0 -3607
rect 33 -3650 66 -3607
rect 0 -3650 33 -3607
rect 99 -3650 132 -3607
rect 165 -3650 198 -3607
rect 198 -3650 231 -3607
rect 231 -3650 264 -3607
rect 297 -3650 330 -3607
rect 330 -3650 363 -3607
rect 363 -3650 396 -3607
rect 429 -3650 462 -3607
rect 396 -3650 429 -3607
rect 495 -3650 528 -3607
rect 561 -3650 594 -3607
rect 528 -3650 561 -3607
rect 627 -3650 660 -3607
rect 693 -3650 726 -3607
rect 726 -3650 759 -3607
rect 759 -3650 792 -3607
rect 825 -3650 858 -3607
rect 792 -3650 825 -3607
rect 891 -3650 924 -3607
rect -53 -3721 -33 -3678
rect -33 -3721 0 -3678
rect 33 -3721 66 -3678
rect 0 -3721 33 -3678
rect 99 -3721 132 -3678
rect 165 -3721 198 -3678
rect 198 -3721 231 -3678
rect 231 -3721 264 -3678
rect 297 -3721 330 -3678
rect 330 -3721 363 -3678
rect 363 -3721 396 -3678
rect 429 -3721 462 -3678
rect 396 -3721 429 -3678
rect 495 -3721 528 -3678
rect 561 -3721 594 -3678
rect 528 -3721 561 -3678
rect 627 -3721 660 -3678
rect 693 -3721 726 -3678
rect 726 -3721 759 -3678
rect 759 -3721 792 -3678
rect 825 -3721 858 -3678
rect 858 -3721 891 -3678
rect 891 -3721 924 -3678
rect -53 -3792 -33 -3749
rect -33 -3792 0 -3749
rect 33 -3792 66 -3749
rect 0 -3792 33 -3749
rect 99 -3792 132 -3749
rect 165 -3792 198 -3749
rect 198 -3792 231 -3749
rect 231 -3792 264 -3749
rect 297 -3792 330 -3749
rect 330 -3792 363 -3749
rect 363 -3792 396 -3749
rect 429 -3792 462 -3749
rect 396 -3792 429 -3749
rect 495 -3792 528 -3749
rect 561 -3792 594 -3749
rect 594 -3792 627 -3749
rect 627 -3792 660 -3749
rect 693 -3792 726 -3749
rect 660 -3792 693 -3749
rect 759 -3792 792 -3749
rect 825 -3792 858 -3749
rect 792 -3792 825 -3749
rect 891 -3792 924 -3749
rect -53 -3863 -33 -3820
rect -33 -3863 0 -3820
rect 33 -3863 66 -3820
rect 0 -3863 33 -3820
rect 99 -3863 132 -3820
rect 165 -3863 198 -3820
rect 198 -3863 231 -3820
rect 231 -3863 264 -3820
rect 297 -3863 330 -3820
rect 330 -3863 363 -3820
rect 363 -3863 396 -3820
rect 429 -3863 462 -3820
rect 396 -3863 429 -3820
rect 495 -3863 528 -3820
rect 561 -3863 594 -3820
rect 594 -3863 627 -3820
rect 627 -3863 660 -3820
rect 693 -3863 726 -3820
rect 660 -3863 693 -3820
rect 759 -3863 792 -3820
rect 825 -3863 858 -3820
rect 858 -3863 891 -3820
rect 891 -3863 924 -3820
rect -53 -3934 -33 -3891
rect -33 -3934 0 -3891
rect 33 -3934 66 -3891
rect 0 -3934 33 -3891
rect 99 -3934 132 -3891
rect 165 -3934 198 -3891
rect 198 -3934 231 -3891
rect 231 -3934 264 -3891
rect 297 -3934 330 -3891
rect 330 -3934 363 -3891
rect 363 -3934 396 -3891
rect 429 -3934 462 -3891
rect 396 -3934 429 -3891
rect 495 -3934 528 -3891
rect 561 -3934 594 -3891
rect 594 -3934 627 -3891
rect 627 -3934 660 -3891
rect 693 -3934 726 -3891
rect 726 -3934 759 -3891
rect 759 -3934 792 -3891
rect 825 -3934 858 -3891
rect 792 -3934 825 -3891
rect 891 -3934 924 -3891
rect -53 -4005 -33 -3962
rect -33 -4005 0 -3962
rect 33 -4005 66 -3962
rect 0 -4005 33 -3962
rect 99 -4005 132 -3962
rect 165 -4005 198 -3962
rect 198 -4005 231 -3962
rect 231 -4005 264 -3962
rect 297 -4005 330 -3962
rect 330 -4005 363 -3962
rect 363 -4005 396 -3962
rect 429 -4005 462 -3962
rect 396 -4005 429 -3962
rect 495 -4005 528 -3962
rect 561 -4005 594 -3962
rect 594 -4005 627 -3962
rect 627 -4005 660 -3962
rect 693 -4005 726 -3962
rect 726 -4005 759 -3962
rect 759 -4005 792 -3962
rect 825 -4005 858 -3962
rect 858 -4005 891 -3962
rect 891 -4005 924 -3962
rect -53 -4076 -33 -4033
rect -33 -4076 0 -4033
rect 33 -4076 66 -4033
rect 0 -4076 33 -4033
rect 99 -4076 132 -4033
rect 165 -4076 198 -4033
rect 198 -4076 231 -4033
rect 231 -4076 264 -4033
rect 297 -4076 330 -4033
rect 330 -4076 363 -4033
rect 363 -4076 396 -4033
rect 429 -4076 462 -4033
rect 462 -4076 495 -4033
rect 495 -4076 528 -4033
rect 561 -4076 594 -4033
rect 528 -4076 561 -4033
rect 627 -4076 660 -4033
rect 693 -4076 726 -4033
rect 660 -4076 693 -4033
rect 759 -4076 792 -4033
rect 825 -4076 858 -4033
rect 792 -4076 825 -4033
rect 891 -4076 924 -4033
rect -53 -4147 -33 -4104
rect -33 -4147 0 -4104
rect 33 -4147 66 -4104
rect 0 -4147 33 -4104
rect 99 -4147 132 -4104
rect 165 -4147 198 -4104
rect 198 -4147 231 -4104
rect 231 -4147 264 -4104
rect 297 -4147 330 -4104
rect 330 -4147 363 -4104
rect 363 -4147 396 -4104
rect 429 -4147 462 -4104
rect 462 -4147 495 -4104
rect 495 -4147 528 -4104
rect 561 -4147 594 -4104
rect 528 -4147 561 -4104
rect 627 -4147 660 -4104
rect 693 -4147 726 -4104
rect 660 -4147 693 -4104
rect 759 -4147 792 -4104
rect 825 -4147 858 -4104
rect 858 -4147 891 -4104
rect 891 -4147 924 -4104
rect -53 -4218 -33 -4175
rect -33 -4218 0 -4175
rect 33 -4218 66 -4175
rect 0 -4218 33 -4175
rect 99 -4218 132 -4175
rect 165 -4218 198 -4175
rect 198 -4218 231 -4175
rect 231 -4218 264 -4175
rect 297 -4218 330 -4175
rect 330 -4218 363 -4175
rect 363 -4218 396 -4175
rect 429 -4218 462 -4175
rect 462 -4218 495 -4175
rect 495 -4218 528 -4175
rect 561 -4218 594 -4175
rect 528 -4218 561 -4175
rect 627 -4218 660 -4175
rect 693 -4218 726 -4175
rect 726 -4218 759 -4175
rect 759 -4218 792 -4175
rect 825 -4218 858 -4175
rect 792 -4218 825 -4175
rect 891 -4218 924 -4175
rect -53 -4289 -33 -4246
rect -33 -4289 0 -4246
rect 33 -4289 66 -4246
rect 0 -4289 33 -4246
rect 99 -4289 132 -4246
rect 165 -4289 198 -4246
rect 198 -4289 231 -4246
rect 231 -4289 264 -4246
rect 297 -4289 330 -4246
rect 330 -4289 363 -4246
rect 363 -4289 396 -4246
rect 429 -4289 462 -4246
rect 462 -4289 495 -4246
rect 495 -4289 528 -4246
rect 561 -4289 594 -4246
rect 528 -4289 561 -4246
rect 627 -4289 660 -4246
rect 693 -4289 726 -4246
rect 726 -4289 759 -4246
rect 759 -4289 792 -4246
rect 825 -4289 858 -4246
rect 858 -4289 891 -4246
rect 891 -4289 924 -4246
rect -53 -4360 -33 -4317
rect -33 -4360 0 -4317
rect 33 -4360 66 -4317
rect 0 -4360 33 -4317
rect 99 -4360 132 -4317
rect 165 -4360 198 -4317
rect 198 -4360 231 -4317
rect 231 -4360 264 -4317
rect 297 -4360 330 -4317
rect 330 -4360 363 -4317
rect 363 -4360 396 -4317
rect 429 -4360 462 -4317
rect 462 -4360 495 -4317
rect 495 -4360 528 -4317
rect 561 -4360 594 -4317
rect 594 -4360 627 -4317
rect 627 -4360 660 -4317
rect 693 -4360 726 -4317
rect 660 -4360 693 -4317
rect 759 -4360 792 -4317
rect 825 -4360 858 -4317
rect 792 -4360 825 -4317
rect 891 -4360 924 -4317
rect -53 -4431 -33 -4388
rect -33 -4431 0 -4388
rect 33 -4431 66 -4388
rect 0 -4431 33 -4388
rect 99 -4431 132 -4388
rect 165 -4431 198 -4388
rect 198 -4431 231 -4388
rect 231 -4431 264 -4388
rect 297 -4431 330 -4388
rect 330 -4431 363 -4388
rect 363 -4431 396 -4388
rect 429 -4431 462 -4388
rect 462 -4431 495 -4388
rect 495 -4431 528 -4388
rect 561 -4431 594 -4388
rect 594 -4431 627 -4388
rect 627 -4431 660 -4388
rect 693 -4431 726 -4388
rect 660 -4431 693 -4388
rect 759 -4431 792 -4388
rect 825 -4431 858 -4388
rect 858 -4431 891 -4388
rect 891 -4431 924 -4388
rect -53 -4502 -33 -4459
rect -33 -4502 0 -4459
rect 33 -4502 66 -4459
rect 0 -4502 33 -4459
rect 99 -4502 132 -4459
rect 165 -4502 198 -4459
rect 198 -4502 231 -4459
rect 231 -4502 264 -4459
rect 297 -4502 330 -4459
rect 330 -4502 363 -4459
rect 363 -4502 396 -4459
rect 429 -4502 462 -4459
rect 462 -4502 495 -4459
rect 495 -4502 528 -4459
rect 561 -4502 594 -4459
rect 594 -4502 627 -4459
rect 627 -4502 660 -4459
rect 693 -4502 726 -4459
rect 726 -4502 759 -4459
rect 759 -4502 792 -4459
rect 825 -4502 858 -4459
rect 792 -4502 825 -4459
rect 891 -4502 924 -4459
rect -53 -4573 -33 -4530
rect -33 -4573 0 -4530
rect 33 -4573 66 -4530
rect 0 -4573 33 -4530
rect 99 -4573 132 -4530
rect 165 -4573 198 -4530
rect 198 -4573 231 -4530
rect 231 -4573 264 -4530
rect 297 -4573 330 -4530
rect 330 -4573 363 -4530
rect 363 -4573 396 -4530
rect 429 -4573 462 -4530
rect 462 -4573 495 -4530
rect 495 -4573 528 -4530
rect 561 -4573 594 -4530
rect 594 -4573 627 -4530
rect 627 -4573 660 -4530
rect 693 -4573 726 -4530
rect 726 -4573 759 -4530
rect 759 -4573 792 -4530
rect 825 -4573 858 -4530
rect 858 -4573 891 -4530
rect 891 -4573 924 -4530
rect -53 -4644 -33 -4601
rect -33 -4644 0 -4601
rect 33 -4644 66 -4601
rect 66 -4644 99 -4601
rect 99 -4644 132 -4601
rect 165 -4644 198 -4601
rect 132 -4644 165 -4601
rect 231 -4644 264 -4601
rect 297 -4644 330 -4601
rect 264 -4644 297 -4601
rect 363 -4644 396 -4601
rect 429 -4644 462 -4601
rect 396 -4644 429 -4601
rect 495 -4644 528 -4601
rect 561 -4644 594 -4601
rect 528 -4644 561 -4601
rect 627 -4644 660 -4601
rect 693 -4644 726 -4601
rect 660 -4644 693 -4601
rect 759 -4644 792 -4601
rect 825 -4644 858 -4601
rect 792 -4644 825 -4601
rect 891 -4644 924 -4601
rect -53 -4715 -33 -4672
rect -33 -4715 0 -4672
rect 33 -4715 66 -4672
rect 66 -4715 99 -4672
rect 99 -4715 132 -4672
rect 165 -4715 198 -4672
rect 132 -4715 165 -4672
rect 231 -4715 264 -4672
rect 297 -4715 330 -4672
rect 264 -4715 297 -4672
rect 363 -4715 396 -4672
rect 429 -4715 462 -4672
rect 396 -4715 429 -4672
rect 495 -4715 528 -4672
rect 561 -4715 594 -4672
rect 528 -4715 561 -4672
rect 627 -4715 660 -4672
rect 693 -4715 726 -4672
rect 660 -4715 693 -4672
rect 759 -4715 792 -4672
rect 825 -4715 858 -4672
rect 858 -4715 891 -4672
rect 891 -4715 924 -4672
rect -53 -4786 -33 -4743
rect -33 -4786 0 -4743
rect 33 -4786 66 -4743
rect 66 -4786 99 -4743
rect 99 -4786 132 -4743
rect 165 -4786 198 -4743
rect 132 -4786 165 -4743
rect 231 -4786 264 -4743
rect 297 -4786 330 -4743
rect 264 -4786 297 -4743
rect 363 -4786 396 -4743
rect 429 -4786 462 -4743
rect 396 -4786 429 -4743
rect 495 -4786 528 -4743
rect 561 -4786 594 -4743
rect 528 -4786 561 -4743
rect 627 -4786 660 -4743
rect 693 -4786 726 -4743
rect 726 -4786 759 -4743
rect 759 -4786 792 -4743
rect 825 -4786 858 -4743
rect 792 -4786 825 -4743
rect 891 -4786 924 -4743
rect -53 -4857 -33 -4814
rect -33 -4857 0 -4814
rect 33 -4857 66 -4814
rect 66 -4857 99 -4814
rect 99 -4857 132 -4814
rect 165 -4857 198 -4814
rect 132 -4857 165 -4814
rect 231 -4857 264 -4814
rect 297 -4857 330 -4814
rect 264 -4857 297 -4814
rect 363 -4857 396 -4814
rect 429 -4857 462 -4814
rect 396 -4857 429 -4814
rect 495 -4857 528 -4814
rect 561 -4857 594 -4814
rect 528 -4857 561 -4814
rect 627 -4857 660 -4814
rect 693 -4857 726 -4814
rect 726 -4857 759 -4814
rect 759 -4857 792 -4814
rect 825 -4857 858 -4814
rect 858 -4857 891 -4814
rect 891 -4857 924 -4814
rect -53 -4928 -33 -4885
rect -33 -4928 0 -4885
rect 33 -4928 66 -4885
rect 66 -4928 99 -4885
rect 99 -4928 132 -4885
rect 165 -4928 198 -4885
rect 132 -4928 165 -4885
rect 231 -4928 264 -4885
rect 297 -4928 330 -4885
rect 264 -4928 297 -4885
rect 363 -4928 396 -4885
rect 429 -4928 462 -4885
rect 396 -4928 429 -4885
rect 495 -4928 528 -4885
rect 561 -4928 594 -4885
rect 594 -4928 627 -4885
rect 627 -4928 660 -4885
rect 693 -4928 726 -4885
rect 660 -4928 693 -4885
rect 759 -4928 792 -4885
rect 825 -4928 858 -4885
rect 792 -4928 825 -4885
rect 891 -4928 924 -4885
rect -53 -4999 -33 -4956
rect -33 -4999 0 -4956
rect 33 -4999 66 -4956
rect 66 -4999 99 -4956
rect 99 -4999 132 -4956
rect 165 -4999 198 -4956
rect 132 -4999 165 -4956
rect 231 -4999 264 -4956
rect 297 -4999 330 -4956
rect 264 -4999 297 -4956
rect 363 -4999 396 -4956
rect 429 -4999 462 -4956
rect 396 -4999 429 -4956
rect 495 -4999 528 -4956
rect 561 -4999 594 -4956
rect 594 -4999 627 -4956
rect 627 -4999 660 -4956
rect 693 -4999 726 -4956
rect 660 -4999 693 -4956
rect 759 -4999 792 -4956
rect 825 -4999 858 -4956
rect 858 -4999 891 -4956
rect 891 -4999 924 -4956
rect -53 -5070 -33 -5027
rect -33 -5070 0 -5027
rect 33 -5070 66 -5027
rect 66 -5070 99 -5027
rect 99 -5070 132 -5027
rect 165 -5070 198 -5027
rect 132 -5070 165 -5027
rect 231 -5070 264 -5027
rect 297 -5070 330 -5027
rect 264 -5070 297 -5027
rect 363 -5070 396 -5027
rect 429 -5070 462 -5027
rect 396 -5070 429 -5027
rect 495 -5070 528 -5027
rect 561 -5070 594 -5027
rect 594 -5070 627 -5027
rect 627 -5070 660 -5027
rect 693 -5070 726 -5027
rect 726 -5070 759 -5027
rect 759 -5070 792 -5027
rect 825 -5070 858 -5027
rect 792 -5070 825 -5027
rect 891 -5070 924 -5027
rect -53 -5141 -33 -5098
rect -33 -5141 0 -5098
rect 33 -5141 66 -5098
rect 66 -5141 99 -5098
rect 99 -5141 132 -5098
rect 165 -5141 198 -5098
rect 132 -5141 165 -5098
rect 231 -5141 264 -5098
rect 297 -5141 330 -5098
rect 264 -5141 297 -5098
rect 363 -5141 396 -5098
rect 429 -5141 462 -5098
rect 396 -5141 429 -5098
rect 495 -5141 528 -5098
rect 561 -5141 594 -5098
rect 594 -5141 627 -5098
rect 627 -5141 660 -5098
rect 693 -5141 726 -5098
rect 726 -5141 759 -5098
rect 759 -5141 792 -5098
rect 825 -5141 858 -5098
rect 858 -5141 891 -5098
rect 891 -5141 924 -5098
rect -53 -5212 -33 -5169
rect -33 -5212 0 -5169
rect 33 -5212 66 -5169
rect 66 -5212 99 -5169
rect 99 -5212 132 -5169
rect 165 -5212 198 -5169
rect 132 -5212 165 -5169
rect 231 -5212 264 -5169
rect 297 -5212 330 -5169
rect 264 -5212 297 -5169
rect 363 -5212 396 -5169
rect 429 -5212 462 -5169
rect 462 -5212 495 -5169
rect 495 -5212 528 -5169
rect 561 -5212 594 -5169
rect 528 -5212 561 -5169
rect 627 -5212 660 -5169
rect 693 -5212 726 -5169
rect 660 -5212 693 -5169
rect 759 -5212 792 -5169
rect 825 -5212 858 -5169
rect 792 -5212 825 -5169
rect 891 -5212 924 -5169
rect -53 -5283 -33 -5240
rect -33 -5283 0 -5240
rect 33 -5283 66 -5240
rect 66 -5283 99 -5240
rect 99 -5283 132 -5240
rect 165 -5283 198 -5240
rect 132 -5283 165 -5240
rect 231 -5283 264 -5240
rect 297 -5283 330 -5240
rect 264 -5283 297 -5240
rect 363 -5283 396 -5240
rect 429 -5283 462 -5240
rect 462 -5283 495 -5240
rect 495 -5283 528 -5240
rect 561 -5283 594 -5240
rect 528 -5283 561 -5240
rect 627 -5283 660 -5240
rect 693 -5283 726 -5240
rect 660 -5283 693 -5240
rect 759 -5283 792 -5240
rect 825 -5283 858 -5240
rect 858 -5283 891 -5240
rect 891 -5283 924 -5240
rect -53 -5354 -33 -5311
rect -33 -5354 0 -5311
rect 33 -5354 66 -5311
rect 66 -5354 99 -5311
rect 99 -5354 132 -5311
rect 165 -5354 198 -5311
rect 132 -5354 165 -5311
rect 231 -5354 264 -5311
rect 297 -5354 330 -5311
rect 264 -5354 297 -5311
rect 363 -5354 396 -5311
rect 429 -5354 462 -5311
rect 462 -5354 495 -5311
rect 495 -5354 528 -5311
rect 561 -5354 594 -5311
rect 528 -5354 561 -5311
rect 627 -5354 660 -5311
rect 693 -5354 726 -5311
rect 726 -5354 759 -5311
rect 759 -5354 792 -5311
rect 825 -5354 858 -5311
rect 792 -5354 825 -5311
rect 891 -5354 924 -5311
rect -53 -5425 -33 -5382
rect -33 -5425 0 -5382
rect 33 -5425 66 -5382
rect 66 -5425 99 -5382
rect 99 -5425 132 -5382
rect 165 -5425 198 -5382
rect 132 -5425 165 -5382
rect 231 -5425 264 -5382
rect 297 -5425 330 -5382
rect 264 -5425 297 -5382
rect 363 -5425 396 -5382
rect 429 -5425 462 -5382
rect 462 -5425 495 -5382
rect 495 -5425 528 -5382
rect 561 -5425 594 -5382
rect 528 -5425 561 -5382
rect 627 -5425 660 -5382
rect 693 -5425 726 -5382
rect 726 -5425 759 -5382
rect 759 -5425 792 -5382
rect 825 -5425 858 -5382
rect 858 -5425 891 -5382
rect 891 -5425 924 -5382
rect -53 -5496 -33 -5453
rect -33 -5496 0 -5453
rect 33 -5496 66 -5453
rect 66 -5496 99 -5453
rect 99 -5496 132 -5453
rect 165 -5496 198 -5453
rect 132 -5496 165 -5453
rect 231 -5496 264 -5453
rect 297 -5496 330 -5453
rect 264 -5496 297 -5453
rect 363 -5496 396 -5453
rect 429 -5496 462 -5453
rect 462 -5496 495 -5453
rect 495 -5496 528 -5453
rect 561 -5496 594 -5453
rect 594 -5496 627 -5453
rect 627 -5496 660 -5453
rect 693 -5496 726 -5453
rect 660 -5496 693 -5453
rect 759 -5496 792 -5453
rect 825 -5496 858 -5453
rect 792 -5496 825 -5453
rect 891 -5496 924 -5453
rect -53 -5567 -33 -5524
rect -33 -5567 0 -5524
rect 33 -5567 66 -5524
rect 66 -5567 99 -5524
rect 99 -5567 132 -5524
rect 165 -5567 198 -5524
rect 132 -5567 165 -5524
rect 231 -5567 264 -5524
rect 297 -5567 330 -5524
rect 264 -5567 297 -5524
rect 363 -5567 396 -5524
rect 429 -5567 462 -5524
rect 462 -5567 495 -5524
rect 495 -5567 528 -5524
rect 561 -5567 594 -5524
rect 594 -5567 627 -5524
rect 627 -5567 660 -5524
rect 693 -5567 726 -5524
rect 660 -5567 693 -5524
rect 759 -5567 792 -5524
rect 825 -5567 858 -5524
rect 858 -5567 891 -5524
rect 891 -5567 924 -5524
rect -53 -5638 -33 -5595
rect -33 -5638 0 -5595
rect 33 -5638 66 -5595
rect 66 -5638 99 -5595
rect 99 -5638 132 -5595
rect 165 -5638 198 -5595
rect 132 -5638 165 -5595
rect 231 -5638 264 -5595
rect 297 -5638 330 -5595
rect 264 -5638 297 -5595
rect 363 -5638 396 -5595
rect 429 -5638 462 -5595
rect 462 -5638 495 -5595
rect 495 -5638 528 -5595
rect 561 -5638 594 -5595
rect 594 -5638 627 -5595
rect 627 -5638 660 -5595
rect 693 -5638 726 -5595
rect 726 -5638 759 -5595
rect 759 -5638 792 -5595
rect 825 -5638 858 -5595
rect 792 -5638 825 -5595
rect 891 -5638 924 -5595
rect -53 -5709 -33 -5666
rect -33 -5709 0 -5666
rect 33 -5709 66 -5666
rect 66 -5709 99 -5666
rect 99 -5709 132 -5666
rect 165 -5709 198 -5666
rect 132 -5709 165 -5666
rect 231 -5709 264 -5666
rect 297 -5709 330 -5666
rect 264 -5709 297 -5666
rect 363 -5709 396 -5666
rect 429 -5709 462 -5666
rect 462 -5709 495 -5666
rect 495 -5709 528 -5666
rect 561 -5709 594 -5666
rect 594 -5709 627 -5666
rect 627 -5709 660 -5666
rect 693 -5709 726 -5666
rect 726 -5709 759 -5666
rect 759 -5709 792 -5666
rect 825 -5709 858 -5666
rect 858 -5709 891 -5666
rect 891 -5709 924 -5666
rect -53 -5780 -33 -5737
rect -33 -5780 0 -5737
rect 33 -5780 66 -5737
rect 66 -5780 99 -5737
rect 99 -5780 132 -5737
rect 165 -5780 198 -5737
rect 132 -5780 165 -5737
rect 231 -5780 264 -5737
rect 297 -5780 330 -5737
rect 330 -5780 363 -5737
rect 363 -5780 396 -5737
rect 429 -5780 462 -5737
rect 396 -5780 429 -5737
rect 495 -5780 528 -5737
rect 561 -5780 594 -5737
rect 528 -5780 561 -5737
rect 627 -5780 660 -5737
rect 693 -5780 726 -5737
rect 660 -5780 693 -5737
rect 759 -5780 792 -5737
rect 825 -5780 858 -5737
rect 792 -5780 825 -5737
rect 891 -5780 924 -5737
rect -53 -5851 -33 -5808
rect -33 -5851 0 -5808
rect 33 -5851 66 -5808
rect 66 -5851 99 -5808
rect 99 -5851 132 -5808
rect 165 -5851 198 -5808
rect 132 -5851 165 -5808
rect 231 -5851 264 -5808
rect 297 -5851 330 -5808
rect 330 -5851 363 -5808
rect 363 -5851 396 -5808
rect 429 -5851 462 -5808
rect 396 -5851 429 -5808
rect 495 -5851 528 -5808
rect 561 -5851 594 -5808
rect 528 -5851 561 -5808
rect 627 -5851 660 -5808
rect 693 -5851 726 -5808
rect 660 -5851 693 -5808
rect 759 -5851 792 -5808
rect 825 -5851 858 -5808
rect 858 -5851 891 -5808
rect 891 -5851 924 -5808
rect -53 -5922 -33 -5879
rect -33 -5922 0 -5879
rect 33 -5922 66 -5879
rect 66 -5922 99 -5879
rect 99 -5922 132 -5879
rect 165 -5922 198 -5879
rect 132 -5922 165 -5879
rect 231 -5922 264 -5879
rect 297 -5922 330 -5879
rect 330 -5922 363 -5879
rect 363 -5922 396 -5879
rect 429 -5922 462 -5879
rect 396 -5922 429 -5879
rect 495 -5922 528 -5879
rect 561 -5922 594 -5879
rect 528 -5922 561 -5879
rect 627 -5922 660 -5879
rect 693 -5922 726 -5879
rect 726 -5922 759 -5879
rect 759 -5922 792 -5879
rect 825 -5922 858 -5879
rect 792 -5922 825 -5879
rect 891 -5922 924 -5879
rect -53 -5993 -33 -5950
rect -33 -5993 0 -5950
rect 33 -5993 66 -5950
rect 66 -5993 99 -5950
rect 99 -5993 132 -5950
rect 165 -5993 198 -5950
rect 132 -5993 165 -5950
rect 231 -5993 264 -5950
rect 297 -5993 330 -5950
rect 330 -5993 363 -5950
rect 363 -5993 396 -5950
rect 429 -5993 462 -5950
rect 396 -5993 429 -5950
rect 495 -5993 528 -5950
rect 561 -5993 594 -5950
rect 528 -5993 561 -5950
rect 627 -5993 660 -5950
rect 693 -5993 726 -5950
rect 726 -5993 759 -5950
rect 759 -5993 792 -5950
rect 825 -5993 858 -5950
rect 858 -5993 891 -5950
rect 891 -5993 924 -5950
rect -53 -6064 -33 -6021
rect -33 -6064 0 -6021
rect 33 -6064 66 -6021
rect 66 -6064 99 -6021
rect 99 -6064 132 -6021
rect 165 -6064 198 -6021
rect 132 -6064 165 -6021
rect 231 -6064 264 -6021
rect 297 -6064 330 -6021
rect 330 -6064 363 -6021
rect 363 -6064 396 -6021
rect 429 -6064 462 -6021
rect 396 -6064 429 -6021
rect 495 -6064 528 -6021
rect 561 -6064 594 -6021
rect 594 -6064 627 -6021
rect 627 -6064 660 -6021
rect 693 -6064 726 -6021
rect 660 -6064 693 -6021
rect 759 -6064 792 -6021
rect 825 -6064 858 -6021
rect 792 -6064 825 -6021
rect 891 -6064 924 -6021
rect -53 -6135 -33 -6092
rect -33 -6135 0 -6092
rect 33 -6135 66 -6092
rect 66 -6135 99 -6092
rect 99 -6135 132 -6092
rect 165 -6135 198 -6092
rect 132 -6135 165 -6092
rect 231 -6135 264 -6092
rect 297 -6135 330 -6092
rect 330 -6135 363 -6092
rect 363 -6135 396 -6092
rect 429 -6135 462 -6092
rect 396 -6135 429 -6092
rect 495 -6135 528 -6092
rect 561 -6135 594 -6092
rect 594 -6135 627 -6092
rect 627 -6135 660 -6092
rect 693 -6135 726 -6092
rect 660 -6135 693 -6092
rect 759 -6135 792 -6092
rect 825 -6135 858 -6092
rect 858 -6135 891 -6092
rect 891 -6135 924 -6092
rect -53 -6206 -33 -6163
rect -33 -6206 0 -6163
rect 33 -6206 66 -6163
rect 66 -6206 99 -6163
rect 99 -6206 132 -6163
rect 165 -6206 198 -6163
rect 132 -6206 165 -6163
rect 231 -6206 264 -6163
rect 297 -6206 330 -6163
rect 330 -6206 363 -6163
rect 363 -6206 396 -6163
rect 429 -6206 462 -6163
rect 396 -6206 429 -6163
rect 495 -6206 528 -6163
rect 561 -6206 594 -6163
rect 594 -6206 627 -6163
rect 627 -6206 660 -6163
rect 693 -6206 726 -6163
rect 726 -6206 759 -6163
rect 759 -6206 792 -6163
rect 825 -6206 858 -6163
rect 792 -6206 825 -6163
rect 891 -6206 924 -6163
rect -53 -6277 -33 -6234
rect -33 -6277 0 -6234
rect 33 -6277 66 -6234
rect 66 -6277 99 -6234
rect 99 -6277 132 -6234
rect 165 -6277 198 -6234
rect 132 -6277 165 -6234
rect 231 -6277 264 -6234
rect 297 -6277 330 -6234
rect 330 -6277 363 -6234
rect 363 -6277 396 -6234
rect 429 -6277 462 -6234
rect 396 -6277 429 -6234
rect 495 -6277 528 -6234
rect 561 -6277 594 -6234
rect 594 -6277 627 -6234
rect 627 -6277 660 -6234
rect 693 -6277 726 -6234
rect 726 -6277 759 -6234
rect 759 -6277 792 -6234
rect 825 -6277 858 -6234
rect 858 -6277 891 -6234
rect 891 -6277 924 -6234
rect -53 -6348 -33 -6305
rect -33 -6348 0 -6305
rect 33 -6348 66 -6305
rect 66 -6348 99 -6305
rect 99 -6348 132 -6305
rect 165 -6348 198 -6305
rect 132 -6348 165 -6305
rect 231 -6348 264 -6305
rect 297 -6348 330 -6305
rect 330 -6348 363 -6305
rect 363 -6348 396 -6305
rect 429 -6348 462 -6305
rect 462 -6348 495 -6305
rect 495 -6348 528 -6305
rect 561 -6348 594 -6305
rect 528 -6348 561 -6305
rect 627 -6348 660 -6305
rect 693 -6348 726 -6305
rect 660 -6348 693 -6305
rect 759 -6348 792 -6305
rect 825 -6348 858 -6305
rect 792 -6348 825 -6305
rect 891 -6348 924 -6305
rect -53 -6419 -33 -6376
rect -33 -6419 0 -6376
rect 33 -6419 66 -6376
rect 66 -6419 99 -6376
rect 99 -6419 132 -6376
rect 165 -6419 198 -6376
rect 132 -6419 165 -6376
rect 231 -6419 264 -6376
rect 297 -6419 330 -6376
rect 330 -6419 363 -6376
rect 363 -6419 396 -6376
rect 429 -6419 462 -6376
rect 462 -6419 495 -6376
rect 495 -6419 528 -6376
rect 561 -6419 594 -6376
rect 528 -6419 561 -6376
rect 627 -6419 660 -6376
rect 693 -6419 726 -6376
rect 660 -6419 693 -6376
rect 759 -6419 792 -6376
rect 825 -6419 858 -6376
rect 858 -6419 891 -6376
rect 891 -6419 924 -6376
rect -53 -6490 -33 -6447
rect -33 -6490 0 -6447
rect 33 -6490 66 -6447
rect 66 -6490 99 -6447
rect 99 -6490 132 -6447
rect 165 -6490 198 -6447
rect 132 -6490 165 -6447
rect 231 -6490 264 -6447
rect 297 -6490 330 -6447
rect 330 -6490 363 -6447
rect 363 -6490 396 -6447
rect 429 -6490 462 -6447
rect 462 -6490 495 -6447
rect 495 -6490 528 -6447
rect 561 -6490 594 -6447
rect 528 -6490 561 -6447
rect 627 -6490 660 -6447
rect 693 -6490 726 -6447
rect 726 -6490 759 -6447
rect 759 -6490 792 -6447
rect 825 -6490 858 -6447
rect 792 -6490 825 -6447
rect 891 -6490 924 -6447
rect -53 -6561 -33 -6518
rect -33 -6561 0 -6518
rect 33 -6561 66 -6518
rect 66 -6561 99 -6518
rect 99 -6561 132 -6518
rect 165 -6561 198 -6518
rect 132 -6561 165 -6518
rect 231 -6561 264 -6518
rect 297 -6561 330 -6518
rect 330 -6561 363 -6518
rect 363 -6561 396 -6518
rect 429 -6561 462 -6518
rect 462 -6561 495 -6518
rect 495 -6561 528 -6518
rect 561 -6561 594 -6518
rect 528 -6561 561 -6518
rect 627 -6561 660 -6518
rect 693 -6561 726 -6518
rect 726 -6561 759 -6518
rect 759 -6561 792 -6518
rect 825 -6561 858 -6518
rect 858 -6561 891 -6518
rect 891 -6561 924 -6518
rect -53 -6632 -33 -6589
rect -33 -6632 0 -6589
rect 33 -6632 66 -6589
rect 66 -6632 99 -6589
rect 99 -6632 132 -6589
rect 165 -6632 198 -6589
rect 132 -6632 165 -6589
rect 231 -6632 264 -6589
rect 297 -6632 330 -6589
rect 330 -6632 363 -6589
rect 363 -6632 396 -6589
rect 429 -6632 462 -6589
rect 462 -6632 495 -6589
rect 495 -6632 528 -6589
rect 561 -6632 594 -6589
rect 594 -6632 627 -6589
rect 627 -6632 660 -6589
rect 693 -6632 726 -6589
rect 660 -6632 693 -6589
rect 759 -6632 792 -6589
rect 825 -6632 858 -6589
rect 792 -6632 825 -6589
rect 891 -6632 924 -6589
rect -53 -6703 -33 -6660
rect -33 -6703 0 -6660
rect 33 -6703 66 -6660
rect 66 -6703 99 -6660
rect 99 -6703 132 -6660
rect 165 -6703 198 -6660
rect 132 -6703 165 -6660
rect 231 -6703 264 -6660
rect 297 -6703 330 -6660
rect 330 -6703 363 -6660
rect 363 -6703 396 -6660
rect 429 -6703 462 -6660
rect 462 -6703 495 -6660
rect 495 -6703 528 -6660
rect 561 -6703 594 -6660
rect 594 -6703 627 -6660
rect 627 -6703 660 -6660
rect 693 -6703 726 -6660
rect 660 -6703 693 -6660
rect 759 -6703 792 -6660
rect 825 -6703 858 -6660
rect 858 -6703 891 -6660
rect 891 -6703 924 -6660
rect -53 -6774 -33 -6731
rect -33 -6774 0 -6731
rect 33 -6774 66 -6731
rect 66 -6774 99 -6731
rect 99 -6774 132 -6731
rect 165 -6774 198 -6731
rect 132 -6774 165 -6731
rect 231 -6774 264 -6731
rect 297 -6774 330 -6731
rect 330 -6774 363 -6731
rect 363 -6774 396 -6731
rect 429 -6774 462 -6731
rect 462 -6774 495 -6731
rect 495 -6774 528 -6731
rect 561 -6774 594 -6731
rect 594 -6774 627 -6731
rect 627 -6774 660 -6731
rect 693 -6774 726 -6731
rect 726 -6774 759 -6731
rect 759 -6774 792 -6731
rect 825 -6774 858 -6731
rect 792 -6774 825 -6731
rect 891 -6774 924 -6731
rect -53 -6845 -33 -6802
rect -33 -6845 0 -6802
rect 33 -6845 66 -6802
rect 66 -6845 99 -6802
rect 99 -6845 132 -6802
rect 165 -6845 198 -6802
rect 132 -6845 165 -6802
rect 231 -6845 264 -6802
rect 297 -6845 330 -6802
rect 330 -6845 363 -6802
rect 363 -6845 396 -6802
rect 429 -6845 462 -6802
rect 462 -6845 495 -6802
rect 495 -6845 528 -6802
rect 561 -6845 594 -6802
rect 594 -6845 627 -6802
rect 627 -6845 660 -6802
rect 693 -6845 726 -6802
rect 726 -6845 759 -6802
rect 759 -6845 792 -6802
rect 825 -6845 858 -6802
rect 858 -6845 891 -6802
rect 891 -6845 924 -6802
rect -53 -6916 -33 -6873
rect -33 -6916 0 -6873
rect 33 -6916 66 -6873
rect 66 -6916 99 -6873
rect 99 -6916 132 -6873
rect 165 -6916 198 -6873
rect 198 -6916 231 -6873
rect 231 -6916 264 -6873
rect 297 -6916 330 -6873
rect 264 -6916 297 -6873
rect 363 -6916 396 -6873
rect 429 -6916 462 -6873
rect 396 -6916 429 -6873
rect 495 -6916 528 -6873
rect 561 -6916 594 -6873
rect 528 -6916 561 -6873
rect 627 -6916 660 -6873
rect 693 -6916 726 -6873
rect 660 -6916 693 -6873
rect 759 -6916 792 -6873
rect 825 -6916 858 -6873
rect 792 -6916 825 -6873
rect 891 -6916 924 -6873
rect -53 -6987 -33 -6944
rect -33 -6987 0 -6944
rect 33 -6987 66 -6944
rect 66 -6987 99 -6944
rect 99 -6987 132 -6944
rect 165 -6987 198 -6944
rect 198 -6987 231 -6944
rect 231 -6987 264 -6944
rect 297 -6987 330 -6944
rect 264 -6987 297 -6944
rect 363 -6987 396 -6944
rect 429 -6987 462 -6944
rect 396 -6987 429 -6944
rect 495 -6987 528 -6944
rect 561 -6987 594 -6944
rect 528 -6987 561 -6944
rect 627 -6987 660 -6944
rect 693 -6987 726 -6944
rect 660 -6987 693 -6944
rect 759 -6987 792 -6944
rect 825 -6987 858 -6944
rect 858 -6987 891 -6944
rect 891 -6987 924 -6944
rect -53 -7058 -33 -7015
rect -33 -7058 0 -7015
rect 33 -7058 66 -7015
rect 66 -7058 99 -7015
rect 99 -7058 132 -7015
rect 165 -7058 198 -7015
rect 198 -7058 231 -7015
rect 231 -7058 264 -7015
rect 297 -7058 330 -7015
rect 264 -7058 297 -7015
rect 363 -7058 396 -7015
rect 429 -7058 462 -7015
rect 396 -7058 429 -7015
rect 495 -7058 528 -7015
rect 561 -7058 594 -7015
rect 528 -7058 561 -7015
rect 627 -7058 660 -7015
rect 693 -7058 726 -7015
rect 726 -7058 759 -7015
rect 759 -7058 792 -7015
rect 825 -7058 858 -7015
rect 792 -7058 825 -7015
rect 891 -7058 924 -7015
rect -53 -7129 -33 -7086
rect -33 -7129 0 -7086
rect 33 -7129 66 -7086
rect 66 -7129 99 -7086
rect 99 -7129 132 -7086
rect 165 -7129 198 -7086
rect 198 -7129 231 -7086
rect 231 -7129 264 -7086
rect 297 -7129 330 -7086
rect 264 -7129 297 -7086
rect 363 -7129 396 -7086
rect 429 -7129 462 -7086
rect 396 -7129 429 -7086
rect 495 -7129 528 -7086
rect 561 -7129 594 -7086
rect 528 -7129 561 -7086
rect 627 -7129 660 -7086
rect 693 -7129 726 -7086
rect 726 -7129 759 -7086
rect 759 -7129 792 -7086
rect 825 -7129 858 -7086
rect 858 -7129 891 -7086
rect 891 -7129 924 -7086
rect -53 -7200 -33 -7157
rect -33 -7200 0 -7157
rect 33 -7200 66 -7157
rect 66 -7200 99 -7157
rect 99 -7200 132 -7157
rect 165 -7200 198 -7157
rect 198 -7200 231 -7157
rect 231 -7200 264 -7157
rect 297 -7200 330 -7157
rect 264 -7200 297 -7157
rect 363 -7200 396 -7157
rect 429 -7200 462 -7157
rect 396 -7200 429 -7157
rect 495 -7200 528 -7157
rect 561 -7200 594 -7157
rect 594 -7200 627 -7157
rect 627 -7200 660 -7157
rect 693 -7200 726 -7157
rect 660 -7200 693 -7157
rect 759 -7200 792 -7157
rect 825 -7200 858 -7157
rect 792 -7200 825 -7157
rect 891 -7200 924 -7157
rect -53 -7271 -33 -7228
rect -33 -7271 0 -7228
rect 33 -7271 66 -7228
rect 66 -7271 99 -7228
rect 99 -7271 132 -7228
rect 165 -7271 198 -7228
rect 198 -7271 231 -7228
rect 231 -7271 264 -7228
rect 297 -7271 330 -7228
rect 264 -7271 297 -7228
rect 363 -7271 396 -7228
rect 429 -7271 462 -7228
rect 396 -7271 429 -7228
rect 495 -7271 528 -7228
rect 561 -7271 594 -7228
rect 594 -7271 627 -7228
rect 627 -7271 660 -7228
rect 693 -7271 726 -7228
rect 660 -7271 693 -7228
rect 759 -7271 792 -7228
rect 825 -7271 858 -7228
rect 858 -7271 891 -7228
rect 891 -7271 924 -7228
rect -53 -7342 -33 -7299
rect -33 -7342 0 -7299
rect 33 -7342 66 -7299
rect 66 -7342 99 -7299
rect 99 -7342 132 -7299
rect 165 -7342 198 -7299
rect 198 -7342 231 -7299
rect 231 -7342 264 -7299
rect 297 -7342 330 -7299
rect 264 -7342 297 -7299
rect 363 -7342 396 -7299
rect 429 -7342 462 -7299
rect 396 -7342 429 -7299
rect 495 -7342 528 -7299
rect 561 -7342 594 -7299
rect 594 -7342 627 -7299
rect 627 -7342 660 -7299
rect 693 -7342 726 -7299
rect 726 -7342 759 -7299
rect 759 -7342 792 -7299
rect 825 -7342 858 -7299
rect 792 -7342 825 -7299
rect 891 -7342 924 -7299
rect -53 -7413 -33 -7370
rect -33 -7413 0 -7370
rect 33 -7413 66 -7370
rect 66 -7413 99 -7370
rect 99 -7413 132 -7370
rect 165 -7413 198 -7370
rect 198 -7413 231 -7370
rect 231 -7413 264 -7370
rect 297 -7413 330 -7370
rect 264 -7413 297 -7370
rect 363 -7413 396 -7370
rect 429 -7413 462 -7370
rect 396 -7413 429 -7370
rect 495 -7413 528 -7370
rect 561 -7413 594 -7370
rect 594 -7413 627 -7370
rect 627 -7413 660 -7370
rect 693 -7413 726 -7370
rect 726 -7413 759 -7370
rect 759 -7413 792 -7370
rect 825 -7413 858 -7370
rect 858 -7413 891 -7370
rect 891 -7413 924 -7370
rect -53 -7484 -33 -7441
rect -33 -7484 0 -7441
rect 33 -7484 66 -7441
rect 66 -7484 99 -7441
rect 99 -7484 132 -7441
rect 165 -7484 198 -7441
rect 198 -7484 231 -7441
rect 231 -7484 264 -7441
rect 297 -7484 330 -7441
rect 264 -7484 297 -7441
rect 363 -7484 396 -7441
rect 429 -7484 462 -7441
rect 462 -7484 495 -7441
rect 495 -7484 528 -7441
rect 561 -7484 594 -7441
rect 528 -7484 561 -7441
rect 627 -7484 660 -7441
rect 693 -7484 726 -7441
rect 660 -7484 693 -7441
rect 759 -7484 792 -7441
rect 825 -7484 858 -7441
rect 792 -7484 825 -7441
rect 891 -7484 924 -7441
rect -53 -7555 -33 -7512
rect -33 -7555 0 -7512
rect 33 -7555 66 -7512
rect 66 -7555 99 -7512
rect 99 -7555 132 -7512
rect 165 -7555 198 -7512
rect 198 -7555 231 -7512
rect 231 -7555 264 -7512
rect 297 -7555 330 -7512
rect 264 -7555 297 -7512
rect 363 -7555 396 -7512
rect 429 -7555 462 -7512
rect 462 -7555 495 -7512
rect 495 -7555 528 -7512
rect 561 -7555 594 -7512
rect 528 -7555 561 -7512
rect 627 -7555 660 -7512
rect 693 -7555 726 -7512
rect 660 -7555 693 -7512
rect 759 -7555 792 -7512
rect 825 -7555 858 -7512
rect 858 -7555 891 -7512
rect 891 -7555 924 -7512
rect -53 -7626 -33 -7583
rect -33 -7626 0 -7583
rect 33 -7626 66 -7583
rect 66 -7626 99 -7583
rect 99 -7626 132 -7583
rect 165 -7626 198 -7583
rect 198 -7626 231 -7583
rect 231 -7626 264 -7583
rect 297 -7626 330 -7583
rect 264 -7626 297 -7583
rect 363 -7626 396 -7583
rect 429 -7626 462 -7583
rect 462 -7626 495 -7583
rect 495 -7626 528 -7583
rect 561 -7626 594 -7583
rect 528 -7626 561 -7583
rect 627 -7626 660 -7583
rect 693 -7626 726 -7583
rect 726 -7626 759 -7583
rect 759 -7626 792 -7583
rect 825 -7626 858 -7583
rect 792 -7626 825 -7583
rect 891 -7626 924 -7583
rect -53 -7697 -33 -7654
rect -33 -7697 0 -7654
rect 33 -7697 66 -7654
rect 66 -7697 99 -7654
rect 99 -7697 132 -7654
rect 165 -7697 198 -7654
rect 198 -7697 231 -7654
rect 231 -7697 264 -7654
rect 297 -7697 330 -7654
rect 264 -7697 297 -7654
rect 363 -7697 396 -7654
rect 429 -7697 462 -7654
rect 462 -7697 495 -7654
rect 495 -7697 528 -7654
rect 561 -7697 594 -7654
rect 528 -7697 561 -7654
rect 627 -7697 660 -7654
rect 693 -7697 726 -7654
rect 726 -7697 759 -7654
rect 759 -7697 792 -7654
rect 825 -7697 858 -7654
rect 858 -7697 891 -7654
rect 891 -7697 924 -7654
rect -53 -7768 -33 -7725
rect -33 -7768 0 -7725
rect 33 -7768 66 -7725
rect 66 -7768 99 -7725
rect 99 -7768 132 -7725
rect 165 -7768 198 -7725
rect 198 -7768 231 -7725
rect 231 -7768 264 -7725
rect 297 -7768 330 -7725
rect 264 -7768 297 -7725
rect 363 -7768 396 -7725
rect 429 -7768 462 -7725
rect 462 -7768 495 -7725
rect 495 -7768 528 -7725
rect 561 -7768 594 -7725
rect 594 -7768 627 -7725
rect 627 -7768 660 -7725
rect 693 -7768 726 -7725
rect 660 -7768 693 -7725
rect 759 -7768 792 -7725
rect 825 -7768 858 -7725
rect 792 -7768 825 -7725
rect 891 -7768 924 -7725
rect -53 -7839 -33 -7796
rect -33 -7839 0 -7796
rect 33 -7839 66 -7796
rect 66 -7839 99 -7796
rect 99 -7839 132 -7796
rect 165 -7839 198 -7796
rect 198 -7839 231 -7796
rect 231 -7839 264 -7796
rect 297 -7839 330 -7796
rect 264 -7839 297 -7796
rect 363 -7839 396 -7796
rect 429 -7839 462 -7796
rect 462 -7839 495 -7796
rect 495 -7839 528 -7796
rect 561 -7839 594 -7796
rect 594 -7839 627 -7796
rect 627 -7839 660 -7796
rect 693 -7839 726 -7796
rect 660 -7839 693 -7796
rect 759 -7839 792 -7796
rect 825 -7839 858 -7796
rect 858 -7839 891 -7796
rect 891 -7839 924 -7796
rect -53 -7910 -33 -7867
rect -33 -7910 0 -7867
rect 33 -7910 66 -7867
rect 66 -7910 99 -7867
rect 99 -7910 132 -7867
rect 165 -7910 198 -7867
rect 198 -7910 231 -7867
rect 231 -7910 264 -7867
rect 297 -7910 330 -7867
rect 264 -7910 297 -7867
rect 363 -7910 396 -7867
rect 429 -7910 462 -7867
rect 462 -7910 495 -7867
rect 495 -7910 528 -7867
rect 561 -7910 594 -7867
rect 594 -7910 627 -7867
rect 627 -7910 660 -7867
rect 693 -7910 726 -7867
rect 726 -7910 759 -7867
rect 759 -7910 792 -7867
rect 825 -7910 858 -7867
rect 792 -7910 825 -7867
rect 891 -7910 924 -7867
rect -53 -7981 -33 -7938
rect -33 -7981 0 -7938
rect 33 -7981 66 -7938
rect 66 -7981 99 -7938
rect 99 -7981 132 -7938
rect 165 -7981 198 -7938
rect 198 -7981 231 -7938
rect 231 -7981 264 -7938
rect 297 -7981 330 -7938
rect 264 -7981 297 -7938
rect 363 -7981 396 -7938
rect 429 -7981 462 -7938
rect 462 -7981 495 -7938
rect 495 -7981 528 -7938
rect 561 -7981 594 -7938
rect 594 -7981 627 -7938
rect 627 -7981 660 -7938
rect 693 -7981 726 -7938
rect 726 -7981 759 -7938
rect 759 -7981 792 -7938
rect 825 -7981 858 -7938
rect 858 -7981 891 -7938
rect 891 -7981 924 -7938
rect -53 -8052 -33 -8009
rect -33 -8052 0 -8009
rect 33 -8052 66 -8009
rect 66 -8052 99 -8009
rect 99 -8052 132 -8009
rect 165 -8052 198 -8009
rect 198 -8052 231 -8009
rect 231 -8052 264 -8009
rect 297 -8052 330 -8009
rect 330 -8052 363 -8009
rect 363 -8052 396 -8009
rect 429 -8052 462 -8009
rect 396 -8052 429 -8009
rect 495 -8052 528 -8009
rect 561 -8052 594 -8009
rect 528 -8052 561 -8009
rect 627 -8052 660 -8009
rect 693 -8052 726 -8009
rect 660 -8052 693 -8009
rect 759 -8052 792 -8009
rect 825 -8052 858 -8009
rect 792 -8052 825 -8009
rect 891 -8052 924 -8009
rect -53 -8123 -33 -8080
rect -33 -8123 0 -8080
rect 33 -8123 66 -8080
rect 66 -8123 99 -8080
rect 99 -8123 132 -8080
rect 165 -8123 198 -8080
rect 198 -8123 231 -8080
rect 231 -8123 264 -8080
rect 297 -8123 330 -8080
rect 330 -8123 363 -8080
rect 363 -8123 396 -8080
rect 429 -8123 462 -8080
rect 396 -8123 429 -8080
rect 495 -8123 528 -8080
rect 561 -8123 594 -8080
rect 528 -8123 561 -8080
rect 627 -8123 660 -8080
rect 693 -8123 726 -8080
rect 660 -8123 693 -8080
rect 759 -8123 792 -8080
rect 825 -8123 858 -8080
rect 858 -8123 891 -8080
rect 891 -8123 924 -8080
rect -53 -8194 -33 -8151
rect -33 -8194 0 -8151
rect 33 -8194 66 -8151
rect 66 -8194 99 -8151
rect 99 -8194 132 -8151
rect 165 -8194 198 -8151
rect 198 -8194 231 -8151
rect 231 -8194 264 -8151
rect 297 -8194 330 -8151
rect 330 -8194 363 -8151
rect 363 -8194 396 -8151
rect 429 -8194 462 -8151
rect 396 -8194 429 -8151
rect 495 -8194 528 -8151
rect 561 -8194 594 -8151
rect 528 -8194 561 -8151
rect 627 -8194 660 -8151
rect 693 -8194 726 -8151
rect 726 -8194 759 -8151
rect 759 -8194 792 -8151
rect 825 -8194 858 -8151
rect 792 -8194 825 -8151
rect 891 -8194 924 -8151
rect -53 -8265 -33 -8222
rect -33 -8265 0 -8222
rect 33 -8265 66 -8222
rect 66 -8265 99 -8222
rect 99 -8265 132 -8222
rect 165 -8265 198 -8222
rect 198 -8265 231 -8222
rect 231 -8265 264 -8222
rect 297 -8265 330 -8222
rect 330 -8265 363 -8222
rect 363 -8265 396 -8222
rect 429 -8265 462 -8222
rect 396 -8265 429 -8222
rect 495 -8265 528 -8222
rect 561 -8265 594 -8222
rect 528 -8265 561 -8222
rect 627 -8265 660 -8222
rect 693 -8265 726 -8222
rect 726 -8265 759 -8222
rect 759 -8265 792 -8222
rect 825 -8265 858 -8222
rect 858 -8265 891 -8222
rect 891 -8265 924 -8222
rect -53 -8336 -33 -8293
rect -33 -8336 0 -8293
rect 33 -8336 66 -8293
rect 66 -8336 99 -8293
rect 99 -8336 132 -8293
rect 165 -8336 198 -8293
rect 198 -8336 231 -8293
rect 231 -8336 264 -8293
rect 297 -8336 330 -8293
rect 330 -8336 363 -8293
rect 363 -8336 396 -8293
rect 429 -8336 462 -8293
rect 396 -8336 429 -8293
rect 495 -8336 528 -8293
rect 561 -8336 594 -8293
rect 594 -8336 627 -8293
rect 627 -8336 660 -8293
rect 693 -8336 726 -8293
rect 660 -8336 693 -8293
rect 759 -8336 792 -8293
rect 825 -8336 858 -8293
rect 792 -8336 825 -8293
rect 891 -8336 924 -8293
rect -53 -8407 -33 -8364
rect -33 -8407 0 -8364
rect 33 -8407 66 -8364
rect 66 -8407 99 -8364
rect 99 -8407 132 -8364
rect 165 -8407 198 -8364
rect 198 -8407 231 -8364
rect 231 -8407 264 -8364
rect 297 -8407 330 -8364
rect 330 -8407 363 -8364
rect 363 -8407 396 -8364
rect 429 -8407 462 -8364
rect 396 -8407 429 -8364
rect 495 -8407 528 -8364
rect 561 -8407 594 -8364
rect 594 -8407 627 -8364
rect 627 -8407 660 -8364
rect 693 -8407 726 -8364
rect 660 -8407 693 -8364
rect 759 -8407 792 -8364
rect 825 -8407 858 -8364
rect 858 -8407 891 -8364
rect 891 -8407 924 -8364
rect -53 -8478 -33 -8435
rect -33 -8478 0 -8435
rect 33 -8478 66 -8435
rect 66 -8478 99 -8435
rect 99 -8478 132 -8435
rect 165 -8478 198 -8435
rect 198 -8478 231 -8435
rect 231 -8478 264 -8435
rect 297 -8478 330 -8435
rect 330 -8478 363 -8435
rect 363 -8478 396 -8435
rect 429 -8478 462 -8435
rect 396 -8478 429 -8435
rect 495 -8478 528 -8435
rect 561 -8478 594 -8435
rect 594 -8478 627 -8435
rect 627 -8478 660 -8435
rect 693 -8478 726 -8435
rect 726 -8478 759 -8435
rect 759 -8478 792 -8435
rect 825 -8478 858 -8435
rect 792 -8478 825 -8435
rect 891 -8478 924 -8435
rect -53 -8549 -33 -8506
rect -33 -8549 0 -8506
rect 33 -8549 66 -8506
rect 66 -8549 99 -8506
rect 99 -8549 132 -8506
rect 165 -8549 198 -8506
rect 198 -8549 231 -8506
rect 231 -8549 264 -8506
rect 297 -8549 330 -8506
rect 330 -8549 363 -8506
rect 363 -8549 396 -8506
rect 429 -8549 462 -8506
rect 396 -8549 429 -8506
rect 495 -8549 528 -8506
rect 561 -8549 594 -8506
rect 594 -8549 627 -8506
rect 627 -8549 660 -8506
rect 693 -8549 726 -8506
rect 726 -8549 759 -8506
rect 759 -8549 792 -8506
rect 825 -8549 858 -8506
rect 858 -8549 891 -8506
rect 891 -8549 924 -8506
rect -53 -8620 -33 -8577
rect -33 -8620 0 -8577
rect 33 -8620 66 -8577
rect 66 -8620 99 -8577
rect 99 -8620 132 -8577
rect 165 -8620 198 -8577
rect 198 -8620 231 -8577
rect 231 -8620 264 -8577
rect 297 -8620 330 -8577
rect 330 -8620 363 -8577
rect 363 -8620 396 -8577
rect 429 -8620 462 -8577
rect 462 -8620 495 -8577
rect 495 -8620 528 -8577
rect 561 -8620 594 -8577
rect 528 -8620 561 -8577
rect 627 -8620 660 -8577
rect 693 -8620 726 -8577
rect 660 -8620 693 -8577
rect 759 -8620 792 -8577
rect 825 -8620 858 -8577
rect 792 -8620 825 -8577
rect 891 -8620 924 -8577
rect -53 -8691 -33 -8648
rect -33 -8691 0 -8648
rect 33 -8691 66 -8648
rect 66 -8691 99 -8648
rect 99 -8691 132 -8648
rect 165 -8691 198 -8648
rect 198 -8691 231 -8648
rect 231 -8691 264 -8648
rect 297 -8691 330 -8648
rect 330 -8691 363 -8648
rect 363 -8691 396 -8648
rect 429 -8691 462 -8648
rect 462 -8691 495 -8648
rect 495 -8691 528 -8648
rect 561 -8691 594 -8648
rect 528 -8691 561 -8648
rect 627 -8691 660 -8648
rect 693 -8691 726 -8648
rect 660 -8691 693 -8648
rect 759 -8691 792 -8648
rect 825 -8691 858 -8648
rect 858 -8691 891 -8648
rect 891 -8691 924 -8648
rect -53 -8762 -33 -8719
rect -33 -8762 0 -8719
rect 33 -8762 66 -8719
rect 66 -8762 99 -8719
rect 99 -8762 132 -8719
rect 165 -8762 198 -8719
rect 198 -8762 231 -8719
rect 231 -8762 264 -8719
rect 297 -8762 330 -8719
rect 330 -8762 363 -8719
rect 363 -8762 396 -8719
rect 429 -8762 462 -8719
rect 462 -8762 495 -8719
rect 495 -8762 528 -8719
rect 561 -8762 594 -8719
rect 528 -8762 561 -8719
rect 627 -8762 660 -8719
rect 693 -8762 726 -8719
rect 726 -8762 759 -8719
rect 759 -8762 792 -8719
rect 825 -8762 858 -8719
rect 792 -8762 825 -8719
rect 891 -8762 924 -8719
rect -53 -8833 -33 -8790
rect -33 -8833 0 -8790
rect 33 -8833 66 -8790
rect 66 -8833 99 -8790
rect 99 -8833 132 -8790
rect 165 -8833 198 -8790
rect 198 -8833 231 -8790
rect 231 -8833 264 -8790
rect 297 -8833 330 -8790
rect 330 -8833 363 -8790
rect 363 -8833 396 -8790
rect 429 -8833 462 -8790
rect 462 -8833 495 -8790
rect 495 -8833 528 -8790
rect 561 -8833 594 -8790
rect 528 -8833 561 -8790
rect 627 -8833 660 -8790
rect 693 -8833 726 -8790
rect 726 -8833 759 -8790
rect 759 -8833 792 -8790
rect 825 -8833 858 -8790
rect 858 -8833 891 -8790
rect 891 -8833 924 -8790
rect -53 -8904 -33 -8861
rect -33 -8904 0 -8861
rect 33 -8904 66 -8861
rect 66 -8904 99 -8861
rect 99 -8904 132 -8861
rect 165 -8904 198 -8861
rect 198 -8904 231 -8861
rect 231 -8904 264 -8861
rect 297 -8904 330 -8861
rect 330 -8904 363 -8861
rect 363 -8904 396 -8861
rect 429 -8904 462 -8861
rect 462 -8904 495 -8861
rect 495 -8904 528 -8861
rect 561 -8904 594 -8861
rect 594 -8904 627 -8861
rect 627 -8904 660 -8861
rect 693 -8904 726 -8861
rect 660 -8904 693 -8861
rect 759 -8904 792 -8861
rect 825 -8904 858 -8861
rect 792 -8904 825 -8861
rect 891 -8904 924 -8861
rect -53 -8975 -33 -8932
rect -33 -8975 0 -8932
rect 33 -8975 66 -8932
rect 66 -8975 99 -8932
rect 99 -8975 132 -8932
rect 165 -8975 198 -8932
rect 198 -8975 231 -8932
rect 231 -8975 264 -8932
rect 297 -8975 330 -8932
rect 330 -8975 363 -8932
rect 363 -8975 396 -8932
rect 429 -8975 462 -8932
rect 462 -8975 495 -8932
rect 495 -8975 528 -8932
rect 561 -8975 594 -8932
rect 594 -8975 627 -8932
rect 627 -8975 660 -8932
rect 693 -8975 726 -8932
rect 660 -8975 693 -8932
rect 759 -8975 792 -8932
rect 825 -8975 858 -8932
rect 858 -8975 891 -8932
rect 891 -8975 924 -8932
rect -53 -9046 -33 -9003
rect -33 -9046 0 -9003
rect 33 -9046 66 -9003
rect 66 -9046 99 -9003
rect 99 -9046 132 -9003
rect 165 -9046 198 -9003
rect 198 -9046 231 -9003
rect 231 -9046 264 -9003
rect 297 -9046 330 -9003
rect 330 -9046 363 -9003
rect 363 -9046 396 -9003
rect 429 -9046 462 -9003
rect 462 -9046 495 -9003
rect 495 -9046 528 -9003
rect 561 -9046 594 -9003
rect 594 -9046 627 -9003
rect 627 -9046 660 -9003
rect 693 -9046 726 -9003
rect 726 -9046 759 -9003
rect 759 -9046 792 -9003
rect 825 -9046 858 -9003
rect 792 -9046 825 -9003
rect 891 -9046 924 -9003
rect -53 -9117 -33 -9074
rect -33 -9117 0 -9074
rect 33 -9117 66 -9074
rect 66 -9117 99 -9074
rect 99 -9117 132 -9074
rect 165 -9117 198 -9074
rect 198 -9117 231 -9074
rect 231 -9117 264 -9074
rect 297 -9117 330 -9074
rect 330 -9117 363 -9074
rect 363 -9117 396 -9074
rect 429 -9117 462 -9074
rect 462 -9117 495 -9074
rect 495 -9117 528 -9074
rect 561 -9117 594 -9074
rect 594 -9117 627 -9074
rect 627 -9117 660 -9074
rect 693 -9117 726 -9074
rect 726 -9117 759 -9074
rect 759 -9117 792 -9074
rect 825 -9117 858 -9074
rect 858 -9117 891 -9074
rect 891 -9117 924 -9074
rect 1022 -100 1055 -57
rect 924 -100 1022 -57
rect 1022 -100 1055 -57
rect 1088 -128 1121 -57
rect 1154 -100 1187 -57
rect 1220 -128 1253 -57
rect 1286 -100 1319 -57
rect 1352 -128 1385 -57
rect 1418 -100 1451 -57
rect 1484 -128 1517 -57
rect 1550 -100 1583 -57
rect 1616 -128 1649 -57
rect 1682 -100 1715 -57
rect 1748 -128 1781 -57
rect 1814 -100 1847 -57
rect 1880 -128 1913 -57
rect 1022 -171 1055 -128
rect 924 -171 1022 -128
rect 1022 -171 1055 -128
rect 1088 -199 1121 -128
rect 1154 -171 1187 -128
rect 1220 -199 1253 -128
rect 1286 -171 1319 -128
rect 1352 -199 1385 -128
rect 1418 -171 1451 -128
rect 1484 -199 1517 -128
rect 1550 -171 1583 -128
rect 1616 -199 1649 -128
rect 1682 -171 1715 -128
rect 1748 -199 1781 -128
rect 1814 -171 1847 -128
rect 1880 -199 1913 -128
rect 1022 -242 1055 -199
rect 924 -242 1022 -199
rect 1022 -242 1055 -199
rect 1088 -270 1121 -199
rect 1154 -242 1187 -199
rect 1220 -270 1253 -199
rect 1286 -242 1319 -199
rect 1352 -270 1385 -199
rect 1418 -242 1451 -199
rect 1484 -270 1517 -199
rect 1550 -242 1583 -199
rect 1616 -270 1649 -199
rect 1682 -242 1715 -199
rect 1748 -270 1781 -199
rect 1814 -242 1847 -199
rect 1880 -270 1913 -199
rect 1022 -313 1055 -270
rect 924 -313 1022 -270
rect 1022 -313 1055 -270
rect 1088 -341 1121 -270
rect 1154 -313 1187 -270
rect 1220 -341 1253 -270
rect 1286 -313 1319 -270
rect 1352 -341 1385 -270
rect 1418 -313 1451 -270
rect 1484 -341 1517 -270
rect 1550 -313 1583 -270
rect 1616 -341 1649 -270
rect 1682 -313 1715 -270
rect 1748 -341 1781 -270
rect 1814 -313 1847 -270
rect 1880 -341 1913 -270
rect 1022 -384 1055 -341
rect 924 -384 1022 -341
rect 1022 -384 1055 -341
rect 1088 -412 1121 -341
rect 1154 -384 1187 -341
rect 1220 -412 1253 -341
rect 1286 -384 1319 -341
rect 1352 -412 1385 -341
rect 1418 -384 1451 -341
rect 1484 -412 1517 -341
rect 1550 -384 1583 -341
rect 1616 -412 1649 -341
rect 1682 -384 1715 -341
rect 1748 -412 1781 -341
rect 1814 -384 1847 -341
rect 1880 -412 1913 -341
rect 1022 -455 1055 -412
rect 924 -455 1022 -412
rect 1022 -455 1055 -412
rect 1088 -483 1121 -412
rect 1154 -455 1187 -412
rect 1220 -483 1253 -412
rect 1286 -455 1319 -412
rect 1352 -483 1385 -412
rect 1418 -455 1451 -412
rect 1484 -483 1517 -412
rect 1550 -455 1583 -412
rect 1616 -483 1649 -412
rect 1682 -455 1715 -412
rect 1748 -483 1781 -412
rect 1814 -455 1847 -412
rect 1880 -483 1913 -412
rect 1022 -526 1055 -483
rect 924 -526 1022 -483
rect 1022 -526 1055 -483
rect 1088 -554 1121 -483
rect 1154 -526 1187 -483
rect 1220 -554 1253 -483
rect 1286 -526 1319 -483
rect 1352 -554 1385 -483
rect 1418 -526 1451 -483
rect 1484 -554 1517 -483
rect 1550 -526 1583 -483
rect 1616 -554 1649 -483
rect 1682 -526 1715 -483
rect 1748 -554 1781 -483
rect 1814 -526 1847 -483
rect 1880 -554 1913 -483
rect 1022 -597 1055 -554
rect 924 -597 1022 -554
rect 1022 -597 1055 -554
rect 1088 -625 1121 -554
rect 1154 -597 1187 -554
rect 1220 -625 1253 -554
rect 1286 -597 1319 -554
rect 1352 -625 1385 -554
rect 1418 -597 1451 -554
rect 1484 -625 1517 -554
rect 1550 -597 1583 -554
rect 1616 -625 1649 -554
rect 1682 -597 1715 -554
rect 1748 -625 1781 -554
rect 1814 -597 1847 -554
rect 1880 -625 1913 -554
rect 1022 -668 1055 -625
rect 924 -668 1022 -625
rect 1022 -668 1055 -625
rect 1088 -696 1121 -625
rect 1154 -668 1187 -625
rect 1220 -696 1253 -625
rect 1286 -668 1319 -625
rect 1352 -696 1385 -625
rect 1418 -668 1451 -625
rect 1484 -696 1517 -625
rect 1550 -668 1583 -625
rect 1616 -696 1649 -625
rect 1682 -668 1715 -625
rect 1748 -696 1781 -625
rect 1814 -668 1847 -625
rect 1880 -696 1913 -625
rect 1022 -739 1055 -696
rect 924 -739 1022 -696
rect 1022 -739 1055 -696
rect 1088 -767 1121 -696
rect 1154 -739 1187 -696
rect 1220 -767 1253 -696
rect 1286 -739 1319 -696
rect 1352 -767 1385 -696
rect 1418 -739 1451 -696
rect 1484 -767 1517 -696
rect 1550 -739 1583 -696
rect 1616 -767 1649 -696
rect 1682 -739 1715 -696
rect 1748 -767 1781 -696
rect 1814 -739 1847 -696
rect 1880 -767 1913 -696
rect 1022 -810 1055 -767
rect 924 -810 1022 -767
rect 1022 -810 1055 -767
rect 1088 -838 1121 -767
rect 1154 -810 1187 -767
rect 1220 -838 1253 -767
rect 1286 -810 1319 -767
rect 1352 -838 1385 -767
rect 1418 -810 1451 -767
rect 1484 -838 1517 -767
rect 1550 -810 1583 -767
rect 1616 -838 1649 -767
rect 1682 -810 1715 -767
rect 1748 -838 1781 -767
rect 1814 -810 1847 -767
rect 1880 -838 1913 -767
rect 1022 -881 1055 -838
rect 924 -881 1022 -838
rect 1022 -881 1055 -838
rect 1088 -909 1121 -838
rect 1154 -881 1187 -838
rect 1220 -909 1253 -838
rect 1286 -881 1319 -838
rect 1352 -909 1385 -838
rect 1418 -881 1451 -838
rect 1484 -909 1517 -838
rect 1550 -881 1583 -838
rect 1616 -909 1649 -838
rect 1682 -881 1715 -838
rect 1748 -909 1781 -838
rect 1814 -881 1847 -838
rect 1880 -909 1913 -838
rect 1022 -952 1055 -909
rect 924 -952 1022 -909
rect 1022 -952 1055 -909
rect 1088 -980 1121 -909
rect 1154 -952 1187 -909
rect 1220 -980 1253 -909
rect 1286 -952 1319 -909
rect 1352 -980 1385 -909
rect 1418 -952 1451 -909
rect 1484 -980 1517 -909
rect 1550 -952 1583 -909
rect 1616 -980 1649 -909
rect 1682 -952 1715 -909
rect 1748 -980 1781 -909
rect 1814 -952 1847 -909
rect 1880 -980 1913 -909
rect 1022 -1023 1055 -980
rect 924 -1023 1022 -980
rect 1022 -1023 1055 -980
rect 1088 -1051 1121 -980
rect 1154 -1023 1187 -980
rect 1220 -1051 1253 -980
rect 1286 -1023 1319 -980
rect 1352 -1051 1385 -980
rect 1418 -1023 1451 -980
rect 1484 -1051 1517 -980
rect 1550 -1023 1583 -980
rect 1616 -1051 1649 -980
rect 1682 -1023 1715 -980
rect 1748 -1051 1781 -980
rect 1814 -1023 1847 -980
rect 1880 -1051 1913 -980
rect 1022 -1094 1055 -1051
rect 924 -1094 1022 -1051
rect 1022 -1094 1055 -1051
rect 1088 -1122 1121 -1051
rect 1154 -1094 1187 -1051
rect 1220 -1122 1253 -1051
rect 1286 -1094 1319 -1051
rect 1352 -1122 1385 -1051
rect 1418 -1094 1451 -1051
rect 1484 -1122 1517 -1051
rect 1550 -1094 1583 -1051
rect 1616 -1122 1649 -1051
rect 1682 -1094 1715 -1051
rect 1748 -1122 1781 -1051
rect 1814 -1094 1847 -1051
rect 1880 -1122 1913 -1051
rect 1022 -1165 1055 -1122
rect 924 -1165 1022 -1122
rect 1022 -1165 1055 -1122
rect 1088 -1193 1121 -1122
rect 1154 -1165 1187 -1122
rect 1220 -1193 1253 -1122
rect 1286 -1165 1319 -1122
rect 1352 -1193 1385 -1122
rect 1418 -1165 1451 -1122
rect 1484 -1193 1517 -1122
rect 1550 -1165 1583 -1122
rect 1616 -1193 1649 -1122
rect 1682 -1165 1715 -1122
rect 1748 -1193 1781 -1122
rect 1814 -1165 1847 -1122
rect 1880 -1193 1913 -1122
rect 1022 -1236 1055 -1193
rect 924 -1236 1022 -1193
rect 1022 -1236 1055 -1193
rect 1088 -1264 1121 -1193
rect 1154 -1236 1187 -1193
rect 1220 -1264 1253 -1193
rect 1286 -1236 1319 -1193
rect 1352 -1264 1385 -1193
rect 1418 -1236 1451 -1193
rect 1484 -1264 1517 -1193
rect 1550 -1236 1583 -1193
rect 1616 -1264 1649 -1193
rect 1682 -1236 1715 -1193
rect 1748 -1264 1781 -1193
rect 1814 -1236 1847 -1193
rect 1880 -1264 1913 -1193
rect 1022 -1307 1055 -1264
rect 924 -1307 1022 -1264
rect 1022 -1307 1055 -1264
rect 1088 -1335 1121 -1264
rect 1154 -1307 1187 -1264
rect 1220 -1335 1253 -1264
rect 1286 -1307 1319 -1264
rect 1352 -1335 1385 -1264
rect 1418 -1307 1451 -1264
rect 1484 -1335 1517 -1264
rect 1550 -1307 1583 -1264
rect 1616 -1335 1649 -1264
rect 1682 -1307 1715 -1264
rect 1748 -1335 1781 -1264
rect 1814 -1307 1847 -1264
rect 1880 -1335 1913 -1264
rect 1022 -1378 1055 -1335
rect 924 -1378 1022 -1335
rect 1022 -1378 1055 -1335
rect 1088 -1406 1121 -1335
rect 1154 -1378 1187 -1335
rect 1220 -1406 1253 -1335
rect 1286 -1378 1319 -1335
rect 1352 -1406 1385 -1335
rect 1418 -1378 1451 -1335
rect 1484 -1406 1517 -1335
rect 1550 -1378 1583 -1335
rect 1616 -1406 1649 -1335
rect 1682 -1378 1715 -1335
rect 1748 -1406 1781 -1335
rect 1814 -1378 1847 -1335
rect 1880 -1406 1913 -1335
rect 1022 -1449 1055 -1406
rect 924 -1449 1022 -1406
rect 1022 -1449 1055 -1406
rect 1088 -1477 1121 -1406
rect 1154 -1449 1187 -1406
rect 1220 -1477 1253 -1406
rect 1286 -1449 1319 -1406
rect 1352 -1477 1385 -1406
rect 1418 -1449 1451 -1406
rect 1484 -1477 1517 -1406
rect 1550 -1449 1583 -1406
rect 1616 -1477 1649 -1406
rect 1682 -1449 1715 -1406
rect 1748 -1477 1781 -1406
rect 1814 -1449 1847 -1406
rect 1880 -1477 1913 -1406
rect 1022 -1520 1055 -1477
rect 924 -1520 1022 -1477
rect 1022 -1520 1055 -1477
rect 1088 -1548 1121 -1477
rect 1154 -1520 1187 -1477
rect 1220 -1548 1253 -1477
rect 1286 -1520 1319 -1477
rect 1352 -1548 1385 -1477
rect 1418 -1520 1451 -1477
rect 1484 -1548 1517 -1477
rect 1550 -1520 1583 -1477
rect 1616 -1548 1649 -1477
rect 1682 -1520 1715 -1477
rect 1748 -1548 1781 -1477
rect 1814 -1520 1847 -1477
rect 1880 -1548 1913 -1477
rect 1022 -1591 1055 -1548
rect 924 -1591 1022 -1548
rect 1022 -1591 1055 -1548
rect 1088 -1619 1121 -1548
rect 1154 -1591 1187 -1548
rect 1220 -1619 1253 -1548
rect 1286 -1591 1319 -1548
rect 1352 -1619 1385 -1548
rect 1418 -1591 1451 -1548
rect 1484 -1619 1517 -1548
rect 1550 -1591 1583 -1548
rect 1616 -1619 1649 -1548
rect 1682 -1591 1715 -1548
rect 1748 -1619 1781 -1548
rect 1814 -1591 1847 -1548
rect 1880 -1619 1913 -1548
rect 1022 -1662 1055 -1619
rect 924 -1662 1022 -1619
rect 1022 -1662 1055 -1619
rect 1088 -1690 1121 -1619
rect 1154 -1662 1187 -1619
rect 1220 -1690 1253 -1619
rect 1286 -1662 1319 -1619
rect 1352 -1690 1385 -1619
rect 1418 -1662 1451 -1619
rect 1484 -1690 1517 -1619
rect 1550 -1662 1583 -1619
rect 1616 -1690 1649 -1619
rect 1682 -1662 1715 -1619
rect 1748 -1690 1781 -1619
rect 1814 -1662 1847 -1619
rect 1880 -1690 1913 -1619
rect 1022 -1733 1055 -1690
rect 924 -1733 1022 -1690
rect 1022 -1733 1055 -1690
rect 1088 -1761 1121 -1690
rect 1154 -1733 1187 -1690
rect 1220 -1761 1253 -1690
rect 1286 -1733 1319 -1690
rect 1352 -1761 1385 -1690
rect 1418 -1733 1451 -1690
rect 1484 -1761 1517 -1690
rect 1550 -1733 1583 -1690
rect 1616 -1761 1649 -1690
rect 1682 -1733 1715 -1690
rect 1748 -1761 1781 -1690
rect 1814 -1733 1847 -1690
rect 1880 -1761 1913 -1690
rect 1022 -1804 1055 -1761
rect 924 -1804 1022 -1761
rect 1022 -1804 1055 -1761
rect 1088 -1832 1121 -1761
rect 1154 -1804 1187 -1761
rect 1220 -1832 1253 -1761
rect 1286 -1804 1319 -1761
rect 1352 -1832 1385 -1761
rect 1418 -1804 1451 -1761
rect 1484 -1832 1517 -1761
rect 1550 -1804 1583 -1761
rect 1616 -1832 1649 -1761
rect 1682 -1804 1715 -1761
rect 1748 -1832 1781 -1761
rect 1814 -1804 1847 -1761
rect 1880 -1832 1913 -1761
rect 1022 -1875 1055 -1832
rect 924 -1875 1022 -1832
rect 1022 -1875 1055 -1832
rect 1088 -1903 1121 -1832
rect 1154 -1875 1187 -1832
rect 1220 -1903 1253 -1832
rect 1286 -1875 1319 -1832
rect 1352 -1903 1385 -1832
rect 1418 -1875 1451 -1832
rect 1484 -1903 1517 -1832
rect 1550 -1875 1583 -1832
rect 1616 -1903 1649 -1832
rect 1682 -1875 1715 -1832
rect 1748 -1903 1781 -1832
rect 1814 -1875 1847 -1832
rect 1880 -1903 1913 -1832
rect 1022 -1946 1055 -1903
rect 924 -1946 1022 -1903
rect 1022 -1946 1055 -1903
rect 1088 -1974 1121 -1903
rect 1154 -1946 1187 -1903
rect 1220 -1974 1253 -1903
rect 1286 -1946 1319 -1903
rect 1352 -1974 1385 -1903
rect 1418 -1946 1451 -1903
rect 1484 -1974 1517 -1903
rect 1550 -1946 1583 -1903
rect 1616 -1974 1649 -1903
rect 1682 -1946 1715 -1903
rect 1748 -1974 1781 -1903
rect 1814 -1946 1847 -1903
rect 1880 -1974 1913 -1903
rect 1022 -2017 1055 -1974
rect 924 -2017 1022 -1974
rect 1022 -2017 1055 -1974
rect 1088 -2045 1121 -1974
rect 1154 -2017 1187 -1974
rect 1220 -2045 1253 -1974
rect 1286 -2017 1319 -1974
rect 1352 -2045 1385 -1974
rect 1418 -2017 1451 -1974
rect 1484 -2045 1517 -1974
rect 1550 -2017 1583 -1974
rect 1616 -2045 1649 -1974
rect 1682 -2017 1715 -1974
rect 1748 -2045 1781 -1974
rect 1814 -2017 1847 -1974
rect 1880 -2045 1913 -1974
rect 1022 -2088 1055 -2045
rect 924 -2088 1022 -2045
rect 1022 -2088 1055 -2045
rect 1088 -2116 1121 -2045
rect 1154 -2088 1187 -2045
rect 1220 -2116 1253 -2045
rect 1286 -2088 1319 -2045
rect 1352 -2116 1385 -2045
rect 1418 -2088 1451 -2045
rect 1484 -2116 1517 -2045
rect 1550 -2088 1583 -2045
rect 1616 -2116 1649 -2045
rect 1682 -2088 1715 -2045
rect 1748 -2116 1781 -2045
rect 1814 -2088 1847 -2045
rect 1880 -2116 1913 -2045
rect 1022 -2159 1055 -2116
rect 924 -2159 1022 -2116
rect 1022 -2159 1055 -2116
rect 1088 -2187 1121 -2116
rect 1154 -2159 1187 -2116
rect 1220 -2187 1253 -2116
rect 1286 -2159 1319 -2116
rect 1352 -2187 1385 -2116
rect 1418 -2159 1451 -2116
rect 1484 -2187 1517 -2116
rect 1550 -2159 1583 -2116
rect 1616 -2187 1649 -2116
rect 1682 -2159 1715 -2116
rect 1748 -2187 1781 -2116
rect 1814 -2159 1847 -2116
rect 1880 -2187 1913 -2116
rect 1022 -2230 1055 -2187
rect 924 -2230 1022 -2187
rect 1022 -2230 1055 -2187
rect 1088 -2258 1121 -2187
rect 1154 -2230 1187 -2187
rect 1220 -2258 1253 -2187
rect 1286 -2230 1319 -2187
rect 1352 -2258 1385 -2187
rect 1418 -2230 1451 -2187
rect 1484 -2258 1517 -2187
rect 1550 -2230 1583 -2187
rect 1616 -2258 1649 -2187
rect 1682 -2230 1715 -2187
rect 1748 -2258 1781 -2187
rect 1814 -2230 1847 -2187
rect 1880 -2258 1913 -2187
rect 1022 -2301 1055 -2258
rect 924 -2301 1022 -2258
rect 1022 -2301 1055 -2258
rect 1088 -2329 1121 -2258
rect 1154 -2301 1187 -2258
rect 1220 -2329 1253 -2258
rect 1286 -2301 1319 -2258
rect 1352 -2329 1385 -2258
rect 1418 -2301 1451 -2258
rect 1484 -2329 1517 -2258
rect 1550 -2301 1583 -2258
rect 1616 -2329 1649 -2258
rect 1682 -2301 1715 -2258
rect 1748 -2329 1781 -2258
rect 1814 -2301 1847 -2258
rect 1880 -2329 1913 -2258
rect 1022 -2372 1055 -2329
rect 924 -2372 1022 -2329
rect 1022 -2372 1055 -2329
rect 1088 -2400 1121 -2329
rect 1154 -2372 1187 -2329
rect 1220 -2400 1253 -2329
rect 1286 -2372 1319 -2329
rect 1352 -2400 1385 -2329
rect 1418 -2372 1451 -2329
rect 1484 -2400 1517 -2329
rect 1550 -2372 1583 -2329
rect 1616 -2400 1649 -2329
rect 1682 -2372 1715 -2329
rect 1748 -2400 1781 -2329
rect 1814 -2372 1847 -2329
rect 1880 -2400 1913 -2329
rect 1022 -2443 1055 -2400
rect 924 -2443 1022 -2400
rect 1022 -2443 1055 -2400
rect 1088 -2471 1121 -2400
rect 1154 -2443 1187 -2400
rect 1220 -2471 1253 -2400
rect 1286 -2443 1319 -2400
rect 1352 -2471 1385 -2400
rect 1418 -2443 1451 -2400
rect 1484 -2471 1517 -2400
rect 1550 -2443 1583 -2400
rect 1616 -2471 1649 -2400
rect 1682 -2443 1715 -2400
rect 1748 -2471 1781 -2400
rect 1814 -2443 1847 -2400
rect 1880 -2471 1913 -2400
rect 1022 -2514 1055 -2471
rect 924 -2514 1022 -2471
rect 1022 -2514 1055 -2471
rect 1088 -2542 1121 -2471
rect 1154 -2514 1187 -2471
rect 1220 -2542 1253 -2471
rect 1286 -2514 1319 -2471
rect 1352 -2542 1385 -2471
rect 1418 -2514 1451 -2471
rect 1484 -2542 1517 -2471
rect 1550 -2514 1583 -2471
rect 1616 -2542 1649 -2471
rect 1682 -2514 1715 -2471
rect 1748 -2542 1781 -2471
rect 1814 -2514 1847 -2471
rect 1880 -2542 1913 -2471
rect 1022 -2585 1055 -2542
rect 924 -2585 1022 -2542
rect 1022 -2585 1055 -2542
rect 1088 -2613 1121 -2542
rect 1154 -2585 1187 -2542
rect 1220 -2613 1253 -2542
rect 1286 -2585 1319 -2542
rect 1352 -2613 1385 -2542
rect 1418 -2585 1451 -2542
rect 1484 -2613 1517 -2542
rect 1550 -2585 1583 -2542
rect 1616 -2613 1649 -2542
rect 1682 -2585 1715 -2542
rect 1748 -2613 1781 -2542
rect 1814 -2585 1847 -2542
rect 1880 -2613 1913 -2542
rect 1022 -2656 1055 -2613
rect 924 -2656 1022 -2613
rect 1022 -2656 1055 -2613
rect 1088 -2684 1121 -2613
rect 1154 -2656 1187 -2613
rect 1220 -2684 1253 -2613
rect 1286 -2656 1319 -2613
rect 1352 -2684 1385 -2613
rect 1418 -2656 1451 -2613
rect 1484 -2684 1517 -2613
rect 1550 -2656 1583 -2613
rect 1616 -2684 1649 -2613
rect 1682 -2656 1715 -2613
rect 1748 -2684 1781 -2613
rect 1814 -2656 1847 -2613
rect 1880 -2684 1913 -2613
rect 1022 -2727 1055 -2684
rect 924 -2727 1022 -2684
rect 1022 -2727 1055 -2684
rect 1088 -2755 1121 -2684
rect 1154 -2727 1187 -2684
rect 1220 -2755 1253 -2684
rect 1286 -2727 1319 -2684
rect 1352 -2755 1385 -2684
rect 1418 -2727 1451 -2684
rect 1484 -2755 1517 -2684
rect 1550 -2727 1583 -2684
rect 1616 -2755 1649 -2684
rect 1682 -2727 1715 -2684
rect 1748 -2755 1781 -2684
rect 1814 -2727 1847 -2684
rect 1880 -2755 1913 -2684
rect 1022 -2798 1055 -2755
rect 924 -2798 1022 -2755
rect 1022 -2798 1055 -2755
rect 1088 -2826 1121 -2755
rect 1154 -2798 1187 -2755
rect 1220 -2826 1253 -2755
rect 1286 -2798 1319 -2755
rect 1352 -2826 1385 -2755
rect 1418 -2798 1451 -2755
rect 1484 -2826 1517 -2755
rect 1550 -2798 1583 -2755
rect 1616 -2826 1649 -2755
rect 1682 -2798 1715 -2755
rect 1748 -2826 1781 -2755
rect 1814 -2798 1847 -2755
rect 1880 -2826 1913 -2755
rect 1022 -2869 1055 -2826
rect 924 -2869 1022 -2826
rect 1022 -2869 1055 -2826
rect 1088 -2897 1121 -2826
rect 1154 -2869 1187 -2826
rect 1220 -2897 1253 -2826
rect 1286 -2869 1319 -2826
rect 1352 -2897 1385 -2826
rect 1418 -2869 1451 -2826
rect 1484 -2897 1517 -2826
rect 1550 -2869 1583 -2826
rect 1616 -2897 1649 -2826
rect 1682 -2869 1715 -2826
rect 1748 -2897 1781 -2826
rect 1814 -2869 1847 -2826
rect 1880 -2897 1913 -2826
rect 1022 -2940 1055 -2897
rect 924 -2940 1022 -2897
rect 1022 -2940 1055 -2897
rect 1088 -2968 1121 -2897
rect 1154 -2940 1187 -2897
rect 1220 -2968 1253 -2897
rect 1286 -2940 1319 -2897
rect 1352 -2968 1385 -2897
rect 1418 -2940 1451 -2897
rect 1484 -2968 1517 -2897
rect 1550 -2940 1583 -2897
rect 1616 -2968 1649 -2897
rect 1682 -2940 1715 -2897
rect 1748 -2968 1781 -2897
rect 1814 -2940 1847 -2897
rect 1880 -2968 1913 -2897
rect 1022 -3011 1055 -2968
rect 924 -3011 1022 -2968
rect 1022 -3011 1055 -2968
rect 1088 -3039 1121 -2968
rect 1154 -3011 1187 -2968
rect 1220 -3039 1253 -2968
rect 1286 -3011 1319 -2968
rect 1352 -3039 1385 -2968
rect 1418 -3011 1451 -2968
rect 1484 -3039 1517 -2968
rect 1550 -3011 1583 -2968
rect 1616 -3039 1649 -2968
rect 1682 -3011 1715 -2968
rect 1748 -3039 1781 -2968
rect 1814 -3011 1847 -2968
rect 1880 -3039 1913 -2968
rect 1022 -3082 1055 -3039
rect 924 -3082 1022 -3039
rect 1022 -3082 1055 -3039
rect 1088 -3110 1121 -3039
rect 1154 -3082 1187 -3039
rect 1220 -3110 1253 -3039
rect 1286 -3082 1319 -3039
rect 1352 -3110 1385 -3039
rect 1418 -3082 1451 -3039
rect 1484 -3110 1517 -3039
rect 1550 -3082 1583 -3039
rect 1616 -3110 1649 -3039
rect 1682 -3082 1715 -3039
rect 1748 -3110 1781 -3039
rect 1814 -3082 1847 -3039
rect 1880 -3110 1913 -3039
rect 1022 -3153 1055 -3110
rect 924 -3153 1022 -3110
rect 1022 -3153 1055 -3110
rect 1088 -3181 1121 -3110
rect 1154 -3153 1187 -3110
rect 1220 -3181 1253 -3110
rect 1286 -3153 1319 -3110
rect 1352 -3181 1385 -3110
rect 1418 -3153 1451 -3110
rect 1484 -3181 1517 -3110
rect 1550 -3153 1583 -3110
rect 1616 -3181 1649 -3110
rect 1682 -3153 1715 -3110
rect 1748 -3181 1781 -3110
rect 1814 -3153 1847 -3110
rect 1880 -3181 1913 -3110
rect 1022 -3224 1055 -3181
rect 924 -3224 1022 -3181
rect 1022 -3224 1055 -3181
rect 1088 -3252 1121 -3181
rect 1154 -3224 1187 -3181
rect 1220 -3252 1253 -3181
rect 1286 -3224 1319 -3181
rect 1352 -3252 1385 -3181
rect 1418 -3224 1451 -3181
rect 1484 -3252 1517 -3181
rect 1550 -3224 1583 -3181
rect 1616 -3252 1649 -3181
rect 1682 -3224 1715 -3181
rect 1748 -3252 1781 -3181
rect 1814 -3224 1847 -3181
rect 1880 -3252 1913 -3181
rect 1022 -3295 1055 -3252
rect 924 -3295 1022 -3252
rect 1022 -3295 1055 -3252
rect 1088 -3323 1121 -3252
rect 1154 -3295 1187 -3252
rect 1220 -3323 1253 -3252
rect 1286 -3295 1319 -3252
rect 1352 -3323 1385 -3252
rect 1418 -3295 1451 -3252
rect 1484 -3323 1517 -3252
rect 1550 -3295 1583 -3252
rect 1616 -3323 1649 -3252
rect 1682 -3295 1715 -3252
rect 1748 -3323 1781 -3252
rect 1814 -3295 1847 -3252
rect 1880 -3323 1913 -3252
rect 1022 -3366 1055 -3323
rect 924 -3366 1022 -3323
rect 1022 -3366 1055 -3323
rect 1088 -3394 1121 -3323
rect 1154 -3366 1187 -3323
rect 1220 -3394 1253 -3323
rect 1286 -3366 1319 -3323
rect 1352 -3394 1385 -3323
rect 1418 -3366 1451 -3323
rect 1484 -3394 1517 -3323
rect 1550 -3366 1583 -3323
rect 1616 -3394 1649 -3323
rect 1682 -3366 1715 -3323
rect 1748 -3394 1781 -3323
rect 1814 -3366 1847 -3323
rect 1880 -3394 1913 -3323
rect 1022 -3437 1055 -3394
rect 924 -3437 1022 -3394
rect 1022 -3437 1055 -3394
rect 1088 -3465 1121 -3394
rect 1154 -3437 1187 -3394
rect 1220 -3465 1253 -3394
rect 1286 -3437 1319 -3394
rect 1352 -3465 1385 -3394
rect 1418 -3437 1451 -3394
rect 1484 -3465 1517 -3394
rect 1550 -3437 1583 -3394
rect 1616 -3465 1649 -3394
rect 1682 -3437 1715 -3394
rect 1748 -3465 1781 -3394
rect 1814 -3437 1847 -3394
rect 1880 -3465 1913 -3394
rect 1022 -3508 1055 -3465
rect 924 -3508 1022 -3465
rect 1022 -3508 1055 -3465
rect 1088 -3536 1121 -3465
rect 1154 -3508 1187 -3465
rect 1220 -3536 1253 -3465
rect 1286 -3508 1319 -3465
rect 1352 -3536 1385 -3465
rect 1418 -3508 1451 -3465
rect 1484 -3536 1517 -3465
rect 1550 -3508 1583 -3465
rect 1616 -3536 1649 -3465
rect 1682 -3508 1715 -3465
rect 1748 -3536 1781 -3465
rect 1814 -3508 1847 -3465
rect 1880 -3536 1913 -3465
rect 1022 -3579 1055 -3536
rect 924 -3579 1022 -3536
rect 1022 -3579 1055 -3536
rect 1088 -3607 1121 -3536
rect 1154 -3579 1187 -3536
rect 1220 -3607 1253 -3536
rect 1286 -3579 1319 -3536
rect 1352 -3607 1385 -3536
rect 1418 -3579 1451 -3536
rect 1484 -3607 1517 -3536
rect 1550 -3579 1583 -3536
rect 1616 -3607 1649 -3536
rect 1682 -3579 1715 -3536
rect 1748 -3607 1781 -3536
rect 1814 -3579 1847 -3536
rect 1880 -3607 1913 -3536
rect 1022 -3650 1055 -3607
rect 924 -3650 1022 -3607
rect 1022 -3650 1055 -3607
rect 1088 -3678 1121 -3607
rect 1154 -3650 1187 -3607
rect 1220 -3678 1253 -3607
rect 1286 -3650 1319 -3607
rect 1352 -3678 1385 -3607
rect 1418 -3650 1451 -3607
rect 1484 -3678 1517 -3607
rect 1550 -3650 1583 -3607
rect 1616 -3678 1649 -3607
rect 1682 -3650 1715 -3607
rect 1748 -3678 1781 -3607
rect 1814 -3650 1847 -3607
rect 1880 -3678 1913 -3607
rect 1022 -3721 1055 -3678
rect 924 -3721 1022 -3678
rect 1022 -3721 1055 -3678
rect 1088 -3749 1121 -3678
rect 1154 -3721 1187 -3678
rect 1220 -3749 1253 -3678
rect 1286 -3721 1319 -3678
rect 1352 -3749 1385 -3678
rect 1418 -3721 1451 -3678
rect 1484 -3749 1517 -3678
rect 1550 -3721 1583 -3678
rect 1616 -3749 1649 -3678
rect 1682 -3721 1715 -3678
rect 1748 -3749 1781 -3678
rect 1814 -3721 1847 -3678
rect 1880 -3749 1913 -3678
rect 1022 -3792 1055 -3749
rect 924 -3792 1022 -3749
rect 1022 -3792 1055 -3749
rect 1088 -3820 1121 -3749
rect 1154 -3792 1187 -3749
rect 1220 -3820 1253 -3749
rect 1286 -3792 1319 -3749
rect 1352 -3820 1385 -3749
rect 1418 -3792 1451 -3749
rect 1484 -3820 1517 -3749
rect 1550 -3792 1583 -3749
rect 1616 -3820 1649 -3749
rect 1682 -3792 1715 -3749
rect 1748 -3820 1781 -3749
rect 1814 -3792 1847 -3749
rect 1880 -3820 1913 -3749
rect 1022 -3863 1055 -3820
rect 924 -3863 1022 -3820
rect 1022 -3863 1055 -3820
rect 1088 -3891 1121 -3820
rect 1154 -3863 1187 -3820
rect 1220 -3891 1253 -3820
rect 1286 -3863 1319 -3820
rect 1352 -3891 1385 -3820
rect 1418 -3863 1451 -3820
rect 1484 -3891 1517 -3820
rect 1550 -3863 1583 -3820
rect 1616 -3891 1649 -3820
rect 1682 -3863 1715 -3820
rect 1748 -3891 1781 -3820
rect 1814 -3863 1847 -3820
rect 1880 -3891 1913 -3820
rect 1022 -3934 1055 -3891
rect 924 -3934 1022 -3891
rect 1022 -3934 1055 -3891
rect 1088 -3962 1121 -3891
rect 1154 -3934 1187 -3891
rect 1220 -3962 1253 -3891
rect 1286 -3934 1319 -3891
rect 1352 -3962 1385 -3891
rect 1418 -3934 1451 -3891
rect 1484 -3962 1517 -3891
rect 1550 -3934 1583 -3891
rect 1616 -3962 1649 -3891
rect 1682 -3934 1715 -3891
rect 1748 -3962 1781 -3891
rect 1814 -3934 1847 -3891
rect 1880 -3962 1913 -3891
rect 1022 -4005 1055 -3962
rect 924 -4005 1022 -3962
rect 1022 -4005 1055 -3962
rect 1088 -4033 1121 -3962
rect 1154 -4005 1187 -3962
rect 1220 -4033 1253 -3962
rect 1286 -4005 1319 -3962
rect 1352 -4033 1385 -3962
rect 1418 -4005 1451 -3962
rect 1484 -4033 1517 -3962
rect 1550 -4005 1583 -3962
rect 1616 -4033 1649 -3962
rect 1682 -4005 1715 -3962
rect 1748 -4033 1781 -3962
rect 1814 -4005 1847 -3962
rect 1880 -4033 1913 -3962
rect 1022 -4076 1055 -4033
rect 924 -4076 1022 -4033
rect 1022 -4076 1055 -4033
rect 1088 -4104 1121 -4033
rect 1154 -4076 1187 -4033
rect 1220 -4104 1253 -4033
rect 1286 -4076 1319 -4033
rect 1352 -4104 1385 -4033
rect 1418 -4076 1451 -4033
rect 1484 -4104 1517 -4033
rect 1550 -4076 1583 -4033
rect 1616 -4104 1649 -4033
rect 1682 -4076 1715 -4033
rect 1748 -4104 1781 -4033
rect 1814 -4076 1847 -4033
rect 1880 -4104 1913 -4033
rect 1022 -4147 1055 -4104
rect 924 -4147 1022 -4104
rect 1022 -4147 1055 -4104
rect 1088 -4175 1121 -4104
rect 1154 -4147 1187 -4104
rect 1220 -4175 1253 -4104
rect 1286 -4147 1319 -4104
rect 1352 -4175 1385 -4104
rect 1418 -4147 1451 -4104
rect 1484 -4175 1517 -4104
rect 1550 -4147 1583 -4104
rect 1616 -4175 1649 -4104
rect 1682 -4147 1715 -4104
rect 1748 -4175 1781 -4104
rect 1814 -4147 1847 -4104
rect 1880 -4175 1913 -4104
rect 1022 -4218 1055 -4175
rect 924 -4218 1022 -4175
rect 1022 -4218 1055 -4175
rect 1088 -4246 1121 -4175
rect 1154 -4218 1187 -4175
rect 1220 -4246 1253 -4175
rect 1286 -4218 1319 -4175
rect 1352 -4246 1385 -4175
rect 1418 -4218 1451 -4175
rect 1484 -4246 1517 -4175
rect 1550 -4218 1583 -4175
rect 1616 -4246 1649 -4175
rect 1682 -4218 1715 -4175
rect 1748 -4246 1781 -4175
rect 1814 -4218 1847 -4175
rect 1880 -4246 1913 -4175
rect 1022 -4289 1055 -4246
rect 924 -4289 1022 -4246
rect 1022 -4289 1055 -4246
rect 1088 -4317 1121 -4246
rect 1154 -4289 1187 -4246
rect 1220 -4317 1253 -4246
rect 1286 -4289 1319 -4246
rect 1352 -4317 1385 -4246
rect 1418 -4289 1451 -4246
rect 1484 -4317 1517 -4246
rect 1550 -4289 1583 -4246
rect 1616 -4317 1649 -4246
rect 1682 -4289 1715 -4246
rect 1748 -4317 1781 -4246
rect 1814 -4289 1847 -4246
rect 1880 -4317 1913 -4246
rect 1022 -4360 1055 -4317
rect 924 -4360 1022 -4317
rect 1022 -4360 1055 -4317
rect 1088 -4388 1121 -4317
rect 1154 -4360 1187 -4317
rect 1220 -4388 1253 -4317
rect 1286 -4360 1319 -4317
rect 1352 -4388 1385 -4317
rect 1418 -4360 1451 -4317
rect 1484 -4388 1517 -4317
rect 1550 -4360 1583 -4317
rect 1616 -4388 1649 -4317
rect 1682 -4360 1715 -4317
rect 1748 -4388 1781 -4317
rect 1814 -4360 1847 -4317
rect 1880 -4388 1913 -4317
rect 1022 -4431 1055 -4388
rect 924 -4431 1022 -4388
rect 1022 -4431 1055 -4388
rect 1088 -4459 1121 -4388
rect 1154 -4431 1187 -4388
rect 1220 -4459 1253 -4388
rect 1286 -4431 1319 -4388
rect 1352 -4459 1385 -4388
rect 1418 -4431 1451 -4388
rect 1484 -4459 1517 -4388
rect 1550 -4431 1583 -4388
rect 1616 -4459 1649 -4388
rect 1682 -4431 1715 -4388
rect 1748 -4459 1781 -4388
rect 1814 -4431 1847 -4388
rect 1880 -4459 1913 -4388
rect 1022 -4502 1055 -4459
rect 924 -4502 1022 -4459
rect 1022 -4502 1055 -4459
rect 1088 -4530 1121 -4459
rect 1154 -4502 1187 -4459
rect 1220 -4530 1253 -4459
rect 1286 -4502 1319 -4459
rect 1352 -4530 1385 -4459
rect 1418 -4502 1451 -4459
rect 1484 -4530 1517 -4459
rect 1550 -4502 1583 -4459
rect 1616 -4530 1649 -4459
rect 1682 -4502 1715 -4459
rect 1748 -4530 1781 -4459
rect 1814 -4502 1847 -4459
rect 1880 -4530 1913 -4459
rect 1022 -4573 1055 -4530
rect 924 -4573 1022 -4530
rect 1022 -4573 1055 -4530
rect 1088 -4601 1121 -4530
rect 1154 -4573 1187 -4530
rect 1220 -4601 1253 -4530
rect 1286 -4573 1319 -4530
rect 1352 -4601 1385 -4530
rect 1418 -4573 1451 -4530
rect 1484 -4601 1517 -4530
rect 1550 -4573 1583 -4530
rect 1616 -4601 1649 -4530
rect 1682 -4573 1715 -4530
rect 1748 -4601 1781 -4530
rect 1814 -4573 1847 -4530
rect 1880 -4601 1913 -4530
rect 1022 -4644 1055 -4601
rect 924 -4644 1022 -4601
rect 1022 -4644 1055 -4601
rect 1088 -4672 1121 -4601
rect 1154 -4644 1187 -4601
rect 1220 -4672 1253 -4601
rect 1286 -4644 1319 -4601
rect 1352 -4672 1385 -4601
rect 1418 -4644 1451 -4601
rect 1484 -4672 1517 -4601
rect 1550 -4644 1583 -4601
rect 1616 -4672 1649 -4601
rect 1682 -4644 1715 -4601
rect 1748 -4672 1781 -4601
rect 1814 -4644 1847 -4601
rect 1946 -4644 1979 -4601
rect 1880 -4672 1913 -4601
rect 1022 -4715 1055 -4672
rect 924 -4715 1022 -4672
rect 1022 -4715 1055 -4672
rect 1088 -4743 1121 -4672
rect 1154 -4715 1187 -4672
rect 1220 -4743 1253 -4672
rect 1286 -4715 1319 -4672
rect 1352 -4743 1385 -4672
rect 1418 -4715 1451 -4672
rect 1484 -4743 1517 -4672
rect 1550 -4715 1583 -4672
rect 1616 -4743 1649 -4672
rect 1682 -4715 1715 -4672
rect 1748 -4743 1781 -4672
rect 1814 -4715 1847 -4672
rect 1946 -4715 1979 -4672
rect 1880 -4743 1913 -4672
rect 1022 -4786 1055 -4743
rect 924 -4786 1022 -4743
rect 1022 -4786 1055 -4743
rect 1088 -4814 1121 -4743
rect 1154 -4786 1187 -4743
rect 1220 -4814 1253 -4743
rect 1286 -4786 1319 -4743
rect 1352 -4814 1385 -4743
rect 1418 -4786 1451 -4743
rect 1484 -4814 1517 -4743
rect 1550 -4786 1583 -4743
rect 1616 -4814 1649 -4743
rect 1682 -4786 1715 -4743
rect 1748 -4814 1781 -4743
rect 1814 -4786 1847 -4743
rect 1946 -4786 1979 -4743
rect 1880 -4814 1913 -4743
rect 1022 -4857 1055 -4814
rect 924 -4857 1022 -4814
rect 1022 -4857 1055 -4814
rect 1088 -4885 1121 -4814
rect 1154 -4857 1187 -4814
rect 1220 -4885 1253 -4814
rect 1286 -4857 1319 -4814
rect 1352 -4885 1385 -4814
rect 1418 -4857 1451 -4814
rect 1484 -4885 1517 -4814
rect 1550 -4857 1583 -4814
rect 1616 -4885 1649 -4814
rect 1682 -4857 1715 -4814
rect 1748 -4885 1781 -4814
rect 1814 -4857 1847 -4814
rect 1946 -4857 1979 -4814
rect 1880 -4885 1913 -4814
rect 1022 -4928 1055 -4885
rect 924 -4928 1022 -4885
rect 1022 -4928 1055 -4885
rect 1088 -4956 1121 -4885
rect 1154 -4928 1187 -4885
rect 1220 -4956 1253 -4885
rect 1286 -4928 1319 -4885
rect 1352 -4956 1385 -4885
rect 1418 -4928 1451 -4885
rect 1484 -4956 1517 -4885
rect 1550 -4928 1583 -4885
rect 1616 -4956 1649 -4885
rect 1682 -4928 1715 -4885
rect 1748 -4956 1781 -4885
rect 1814 -4928 1847 -4885
rect 1946 -4928 1979 -4885
rect 1880 -4956 1913 -4885
rect 1022 -4999 1055 -4956
rect 924 -4999 1022 -4956
rect 1022 -4999 1055 -4956
rect 1088 -5027 1121 -4956
rect 1154 -4999 1187 -4956
rect 1220 -5027 1253 -4956
rect 1286 -4999 1319 -4956
rect 1352 -5027 1385 -4956
rect 1418 -4999 1451 -4956
rect 1484 -5027 1517 -4956
rect 1550 -4999 1583 -4956
rect 1616 -5027 1649 -4956
rect 1682 -4999 1715 -4956
rect 1748 -5027 1781 -4956
rect 1814 -4999 1847 -4956
rect 1946 -4999 1979 -4956
rect 1880 -5027 1913 -4956
rect 1022 -5070 1055 -5027
rect 924 -5070 1022 -5027
rect 1022 -5070 1055 -5027
rect 1088 -5098 1121 -5027
rect 1154 -5070 1187 -5027
rect 1220 -5098 1253 -5027
rect 1286 -5070 1319 -5027
rect 1352 -5098 1385 -5027
rect 1418 -5070 1451 -5027
rect 1484 -5098 1517 -5027
rect 1550 -5070 1583 -5027
rect 1616 -5098 1649 -5027
rect 1682 -5070 1715 -5027
rect 1748 -5098 1781 -5027
rect 1814 -5070 1847 -5027
rect 1946 -5070 1979 -5027
rect 1880 -5098 1913 -5027
rect 1022 -5141 1055 -5098
rect 924 -5141 1022 -5098
rect 1022 -5141 1055 -5098
rect 1088 -5169 1121 -5098
rect 1154 -5141 1187 -5098
rect 1220 -5169 1253 -5098
rect 1286 -5141 1319 -5098
rect 1352 -5169 1385 -5098
rect 1418 -5141 1451 -5098
rect 1484 -5169 1517 -5098
rect 1550 -5141 1583 -5098
rect 1616 -5169 1649 -5098
rect 1682 -5141 1715 -5098
rect 1748 -5169 1781 -5098
rect 1814 -5141 1847 -5098
rect 1946 -5141 1979 -5098
rect 1880 -5169 1913 -5098
rect 1022 -5212 1055 -5169
rect 924 -5212 1022 -5169
rect 1022 -5212 1055 -5169
rect 1088 -5240 1121 -5169
rect 1154 -5212 1187 -5169
rect 1220 -5240 1253 -5169
rect 1286 -5212 1319 -5169
rect 1352 -5240 1385 -5169
rect 1418 -5212 1451 -5169
rect 1484 -5240 1517 -5169
rect 1550 -5212 1583 -5169
rect 1616 -5240 1649 -5169
rect 1682 -5212 1715 -5169
rect 1748 -5240 1781 -5169
rect 1814 -5212 1847 -5169
rect 1946 -5212 1979 -5169
rect 1880 -5240 1913 -5169
rect 1022 -5283 1055 -5240
rect 924 -5283 1022 -5240
rect 1022 -5283 1055 -5240
rect 1088 -5311 1121 -5240
rect 1154 -5283 1187 -5240
rect 1220 -5311 1253 -5240
rect 1286 -5283 1319 -5240
rect 1352 -5311 1385 -5240
rect 1418 -5283 1451 -5240
rect 1484 -5311 1517 -5240
rect 1550 -5283 1583 -5240
rect 1616 -5311 1649 -5240
rect 1682 -5283 1715 -5240
rect 1748 -5311 1781 -5240
rect 1814 -5283 1847 -5240
rect 1946 -5283 1979 -5240
rect 1880 -5311 1913 -5240
rect 1022 -5354 1055 -5311
rect 924 -5354 1022 -5311
rect 1022 -5354 1055 -5311
rect 1088 -5382 1121 -5311
rect 1154 -5354 1187 -5311
rect 1220 -5382 1253 -5311
rect 1286 -5354 1319 -5311
rect 1352 -5382 1385 -5311
rect 1418 -5354 1451 -5311
rect 1484 -5382 1517 -5311
rect 1550 -5354 1583 -5311
rect 1616 -5382 1649 -5311
rect 1682 -5354 1715 -5311
rect 1748 -5382 1781 -5311
rect 1814 -5354 1847 -5311
rect 1946 -5354 1979 -5311
rect 1880 -5382 1913 -5311
rect 1022 -5425 1055 -5382
rect 924 -5425 1022 -5382
rect 1022 -5425 1055 -5382
rect 1088 -5453 1121 -5382
rect 1154 -5425 1187 -5382
rect 1220 -5453 1253 -5382
rect 1286 -5425 1319 -5382
rect 1352 -5453 1385 -5382
rect 1418 -5425 1451 -5382
rect 1484 -5453 1517 -5382
rect 1550 -5425 1583 -5382
rect 1616 -5453 1649 -5382
rect 1682 -5425 1715 -5382
rect 1748 -5453 1781 -5382
rect 1814 -5425 1847 -5382
rect 1946 -5425 1979 -5382
rect 1880 -5453 1913 -5382
rect 1022 -5496 1055 -5453
rect 924 -5496 1022 -5453
rect 1022 -5496 1055 -5453
rect 1088 -5524 1121 -5453
rect 1154 -5496 1187 -5453
rect 1220 -5524 1253 -5453
rect 1286 -5496 1319 -5453
rect 1352 -5524 1385 -5453
rect 1418 -5496 1451 -5453
rect 1484 -5524 1517 -5453
rect 1550 -5496 1583 -5453
rect 1616 -5524 1649 -5453
rect 1682 -5496 1715 -5453
rect 1748 -5524 1781 -5453
rect 1814 -5496 1847 -5453
rect 1946 -5496 1979 -5453
rect 1880 -5524 1913 -5453
rect 1022 -5567 1055 -5524
rect 924 -5567 1022 -5524
rect 1022 -5567 1055 -5524
rect 1088 -5595 1121 -5524
rect 1154 -5567 1187 -5524
rect 1220 -5595 1253 -5524
rect 1286 -5567 1319 -5524
rect 1352 -5595 1385 -5524
rect 1418 -5567 1451 -5524
rect 1484 -5595 1517 -5524
rect 1550 -5567 1583 -5524
rect 1616 -5595 1649 -5524
rect 1682 -5567 1715 -5524
rect 1748 -5595 1781 -5524
rect 1814 -5567 1847 -5524
rect 1946 -5567 1979 -5524
rect 1880 -5595 1913 -5524
rect 1022 -5638 1055 -5595
rect 924 -5638 1022 -5595
rect 1022 -5638 1055 -5595
rect 1088 -5666 1121 -5595
rect 1154 -5638 1187 -5595
rect 1220 -5666 1253 -5595
rect 1286 -5638 1319 -5595
rect 1352 -5666 1385 -5595
rect 1418 -5638 1451 -5595
rect 1484 -5666 1517 -5595
rect 1550 -5638 1583 -5595
rect 1616 -5666 1649 -5595
rect 1682 -5638 1715 -5595
rect 1748 -5666 1781 -5595
rect 1814 -5638 1847 -5595
rect 1946 -5638 1979 -5595
rect 1880 -5666 1913 -5595
rect 1022 -5709 1055 -5666
rect 924 -5709 1022 -5666
rect 1022 -5709 1055 -5666
rect 1088 -5737 1121 -5666
rect 1154 -5709 1187 -5666
rect 1220 -5737 1253 -5666
rect 1286 -5709 1319 -5666
rect 1352 -5737 1385 -5666
rect 1418 -5709 1451 -5666
rect 1484 -5737 1517 -5666
rect 1550 -5709 1583 -5666
rect 1616 -5737 1649 -5666
rect 1682 -5709 1715 -5666
rect 1748 -5737 1781 -5666
rect 1814 -5709 1847 -5666
rect 1946 -5709 1979 -5666
rect 1880 -5737 1913 -5666
rect 1022 -5780 1055 -5737
rect 924 -5780 1022 -5737
rect 1022 -5780 1055 -5737
rect 1088 -5808 1121 -5737
rect 1154 -5780 1187 -5737
rect 1220 -5808 1253 -5737
rect 1286 -5780 1319 -5737
rect 1352 -5808 1385 -5737
rect 1418 -5780 1451 -5737
rect 1484 -5808 1517 -5737
rect 1550 -5780 1583 -5737
rect 1616 -5808 1649 -5737
rect 1682 -5780 1715 -5737
rect 1748 -5808 1781 -5737
rect 1814 -5780 1847 -5737
rect 1946 -5780 1979 -5737
rect 1880 -5808 1913 -5737
rect 1022 -5851 1055 -5808
rect 924 -5851 1022 -5808
rect 1022 -5851 1055 -5808
rect 1088 -5879 1121 -5808
rect 1154 -5851 1187 -5808
rect 1220 -5879 1253 -5808
rect 1286 -5851 1319 -5808
rect 1352 -5879 1385 -5808
rect 1418 -5851 1451 -5808
rect 1484 -5879 1517 -5808
rect 1550 -5851 1583 -5808
rect 1616 -5879 1649 -5808
rect 1682 -5851 1715 -5808
rect 1748 -5879 1781 -5808
rect 1814 -5851 1847 -5808
rect 1946 -5851 1979 -5808
rect 1880 -5879 1913 -5808
rect 1022 -5922 1055 -5879
rect 924 -5922 1022 -5879
rect 1022 -5922 1055 -5879
rect 1088 -5950 1121 -5879
rect 1154 -5922 1187 -5879
rect 1220 -5950 1253 -5879
rect 1286 -5922 1319 -5879
rect 1352 -5950 1385 -5879
rect 1418 -5922 1451 -5879
rect 1484 -5950 1517 -5879
rect 1550 -5922 1583 -5879
rect 1616 -5950 1649 -5879
rect 1682 -5922 1715 -5879
rect 1748 -5950 1781 -5879
rect 1814 -5922 1847 -5879
rect 1946 -5922 1979 -5879
rect 1880 -5950 1913 -5879
rect 1022 -5993 1055 -5950
rect 924 -5993 1022 -5950
rect 1022 -5993 1055 -5950
rect 1088 -6021 1121 -5950
rect 1154 -5993 1187 -5950
rect 1220 -6021 1253 -5950
rect 1286 -5993 1319 -5950
rect 1352 -6021 1385 -5950
rect 1418 -5993 1451 -5950
rect 1484 -6021 1517 -5950
rect 1550 -5993 1583 -5950
rect 1616 -6021 1649 -5950
rect 1682 -5993 1715 -5950
rect 1748 -6021 1781 -5950
rect 1814 -5993 1847 -5950
rect 1946 -5993 1979 -5950
rect 1880 -6021 1913 -5950
rect 1022 -6064 1055 -6021
rect 924 -6064 1022 -6021
rect 1022 -6064 1055 -6021
rect 1088 -6092 1121 -6021
rect 1154 -6064 1187 -6021
rect 1220 -6092 1253 -6021
rect 1286 -6064 1319 -6021
rect 1352 -6092 1385 -6021
rect 1418 -6064 1451 -6021
rect 1484 -6092 1517 -6021
rect 1550 -6064 1583 -6021
rect 1616 -6092 1649 -6021
rect 1682 -6064 1715 -6021
rect 1748 -6092 1781 -6021
rect 1814 -6064 1847 -6021
rect 1946 -6064 1979 -6021
rect 1880 -6092 1913 -6021
rect 1022 -6135 1055 -6092
rect 924 -6135 1022 -6092
rect 1022 -6135 1055 -6092
rect 1088 -6163 1121 -6092
rect 1154 -6135 1187 -6092
rect 1220 -6163 1253 -6092
rect 1286 -6135 1319 -6092
rect 1352 -6163 1385 -6092
rect 1418 -6135 1451 -6092
rect 1484 -6163 1517 -6092
rect 1550 -6135 1583 -6092
rect 1616 -6163 1649 -6092
rect 1682 -6135 1715 -6092
rect 1748 -6163 1781 -6092
rect 1814 -6135 1847 -6092
rect 1946 -6135 1979 -6092
rect 1880 -6163 1913 -6092
rect 1022 -6206 1055 -6163
rect 924 -6206 1022 -6163
rect 1022 -6206 1055 -6163
rect 1088 -6234 1121 -6163
rect 1154 -6206 1187 -6163
rect 1220 -6234 1253 -6163
rect 1286 -6206 1319 -6163
rect 1352 -6234 1385 -6163
rect 1418 -6206 1451 -6163
rect 1484 -6234 1517 -6163
rect 1550 -6206 1583 -6163
rect 1616 -6234 1649 -6163
rect 1682 -6206 1715 -6163
rect 1748 -6234 1781 -6163
rect 1814 -6206 1847 -6163
rect 1946 -6206 1979 -6163
rect 1880 -6234 1913 -6163
rect 1022 -6277 1055 -6234
rect 924 -6277 1022 -6234
rect 1022 -6277 1055 -6234
rect 1088 -6305 1121 -6234
rect 1154 -6277 1187 -6234
rect 1220 -6305 1253 -6234
rect 1286 -6277 1319 -6234
rect 1352 -6305 1385 -6234
rect 1418 -6277 1451 -6234
rect 1484 -6305 1517 -6234
rect 1550 -6277 1583 -6234
rect 1616 -6305 1649 -6234
rect 1682 -6277 1715 -6234
rect 1748 -6305 1781 -6234
rect 1814 -6277 1847 -6234
rect 1946 -6277 1979 -6234
rect 1880 -6305 1913 -6234
rect 1022 -6348 1055 -6305
rect 924 -6348 1022 -6305
rect 1022 -6348 1055 -6305
rect 1088 -6376 1121 -6305
rect 1154 -6348 1187 -6305
rect 1220 -6376 1253 -6305
rect 1286 -6348 1319 -6305
rect 1352 -6376 1385 -6305
rect 1418 -6348 1451 -6305
rect 1484 -6376 1517 -6305
rect 1550 -6348 1583 -6305
rect 1616 -6376 1649 -6305
rect 1682 -6348 1715 -6305
rect 1748 -6376 1781 -6305
rect 1814 -6348 1847 -6305
rect 1946 -6348 1979 -6305
rect 1880 -6376 1913 -6305
rect 1022 -6419 1055 -6376
rect 924 -6419 1022 -6376
rect 1022 -6419 1055 -6376
rect 1088 -6447 1121 -6376
rect 1154 -6419 1187 -6376
rect 1220 -6447 1253 -6376
rect 1286 -6419 1319 -6376
rect 1352 -6447 1385 -6376
rect 1418 -6419 1451 -6376
rect 1484 -6447 1517 -6376
rect 1550 -6419 1583 -6376
rect 1616 -6447 1649 -6376
rect 1682 -6419 1715 -6376
rect 1748 -6447 1781 -6376
rect 1814 -6419 1847 -6376
rect 1946 -6419 1979 -6376
rect 1880 -6447 1913 -6376
rect 1022 -6490 1055 -6447
rect 924 -6490 1022 -6447
rect 1022 -6490 1055 -6447
rect 1088 -6518 1121 -6447
rect 1154 -6490 1187 -6447
rect 1220 -6518 1253 -6447
rect 1286 -6490 1319 -6447
rect 1352 -6518 1385 -6447
rect 1418 -6490 1451 -6447
rect 1484 -6518 1517 -6447
rect 1550 -6490 1583 -6447
rect 1616 -6518 1649 -6447
rect 1682 -6490 1715 -6447
rect 1748 -6518 1781 -6447
rect 1814 -6490 1847 -6447
rect 1946 -6490 1979 -6447
rect 1880 -6518 1913 -6447
rect 1022 -6561 1055 -6518
rect 924 -6561 1022 -6518
rect 1022 -6561 1055 -6518
rect 1088 -6589 1121 -6518
rect 1154 -6561 1187 -6518
rect 1220 -6589 1253 -6518
rect 1286 -6561 1319 -6518
rect 1352 -6589 1385 -6518
rect 1418 -6561 1451 -6518
rect 1484 -6589 1517 -6518
rect 1550 -6561 1583 -6518
rect 1616 -6589 1649 -6518
rect 1682 -6561 1715 -6518
rect 1748 -6589 1781 -6518
rect 1814 -6561 1847 -6518
rect 1946 -6561 1979 -6518
rect 1880 -6589 1913 -6518
rect 1022 -6632 1055 -6589
rect 924 -6632 1022 -6589
rect 1022 -6632 1055 -6589
rect 1088 -6660 1121 -6589
rect 1154 -6632 1187 -6589
rect 1220 -6660 1253 -6589
rect 1286 -6632 1319 -6589
rect 1352 -6660 1385 -6589
rect 1418 -6632 1451 -6589
rect 1484 -6660 1517 -6589
rect 1550 -6632 1583 -6589
rect 1616 -6660 1649 -6589
rect 1682 -6632 1715 -6589
rect 1748 -6660 1781 -6589
rect 1814 -6632 1847 -6589
rect 1946 -6632 1979 -6589
rect 1880 -6660 1913 -6589
rect 1022 -6703 1055 -6660
rect 924 -6703 1022 -6660
rect 1022 -6703 1055 -6660
rect 1088 -6731 1121 -6660
rect 1154 -6703 1187 -6660
rect 1220 -6731 1253 -6660
rect 1286 -6703 1319 -6660
rect 1352 -6731 1385 -6660
rect 1418 -6703 1451 -6660
rect 1484 -6731 1517 -6660
rect 1550 -6703 1583 -6660
rect 1616 -6731 1649 -6660
rect 1682 -6703 1715 -6660
rect 1748 -6731 1781 -6660
rect 1814 -6703 1847 -6660
rect 1946 -6703 1979 -6660
rect 1880 -6731 1913 -6660
rect 1022 -6774 1055 -6731
rect 924 -6774 1022 -6731
rect 1022 -6774 1055 -6731
rect 1088 -6802 1121 -6731
rect 1154 -6774 1187 -6731
rect 1220 -6802 1253 -6731
rect 1286 -6774 1319 -6731
rect 1352 -6802 1385 -6731
rect 1418 -6774 1451 -6731
rect 1484 -6802 1517 -6731
rect 1550 -6774 1583 -6731
rect 1616 -6802 1649 -6731
rect 1682 -6774 1715 -6731
rect 1748 -6802 1781 -6731
rect 1814 -6774 1847 -6731
rect 1946 -6774 1979 -6731
rect 1880 -6802 1913 -6731
rect 1022 -6845 1055 -6802
rect 924 -6845 1022 -6802
rect 1022 -6845 1055 -6802
rect 1088 -6873 1121 -6802
rect 1154 -6845 1187 -6802
rect 1220 -6873 1253 -6802
rect 1286 -6845 1319 -6802
rect 1352 -6873 1385 -6802
rect 1418 -6845 1451 -6802
rect 1484 -6873 1517 -6802
rect 1550 -6845 1583 -6802
rect 1616 -6873 1649 -6802
rect 1682 -6845 1715 -6802
rect 1748 -6873 1781 -6802
rect 1814 -6845 1847 -6802
rect 1946 -6845 1979 -6802
rect 1880 -6873 1913 -6802
rect 1022 -6916 1055 -6873
rect 924 -6916 1022 -6873
rect 1022 -6916 1055 -6873
rect 1088 -6944 1121 -6873
rect 1154 -6916 1187 -6873
rect 1220 -6944 1253 -6873
rect 1286 -6916 1319 -6873
rect 1352 -6944 1385 -6873
rect 1418 -6916 1451 -6873
rect 1484 -6944 1517 -6873
rect 1550 -6916 1583 -6873
rect 1616 -6944 1649 -6873
rect 1682 -6916 1715 -6873
rect 1748 -6944 1781 -6873
rect 1814 -6916 1847 -6873
rect 1946 -6916 1979 -6873
rect 1880 -6944 1913 -6873
rect 1022 -6987 1055 -6944
rect 924 -6987 1022 -6944
rect 1022 -6987 1055 -6944
rect 1088 -7015 1121 -6944
rect 1154 -6987 1187 -6944
rect 1220 -7015 1253 -6944
rect 1286 -6987 1319 -6944
rect 1352 -7015 1385 -6944
rect 1418 -6987 1451 -6944
rect 1484 -7015 1517 -6944
rect 1550 -6987 1583 -6944
rect 1616 -7015 1649 -6944
rect 1682 -6987 1715 -6944
rect 1748 -7015 1781 -6944
rect 1814 -6987 1847 -6944
rect 1946 -6987 1979 -6944
rect 1880 -7015 1913 -6944
rect 1022 -7058 1055 -7015
rect 924 -7058 1022 -7015
rect 1022 -7058 1055 -7015
rect 1088 -7086 1121 -7015
rect 1154 -7058 1187 -7015
rect 1220 -7086 1253 -7015
rect 1286 -7058 1319 -7015
rect 1352 -7086 1385 -7015
rect 1418 -7058 1451 -7015
rect 1484 -7086 1517 -7015
rect 1550 -7058 1583 -7015
rect 1616 -7086 1649 -7015
rect 1682 -7058 1715 -7015
rect 1748 -7086 1781 -7015
rect 1814 -7058 1847 -7015
rect 1946 -7058 1979 -7015
rect 1880 -7086 1913 -7015
rect 1022 -7129 1055 -7086
rect 924 -7129 1022 -7086
rect 1022 -7129 1055 -7086
rect 1088 -7157 1121 -7086
rect 1154 -7129 1187 -7086
rect 1220 -7157 1253 -7086
rect 1286 -7129 1319 -7086
rect 1352 -7157 1385 -7086
rect 1418 -7129 1451 -7086
rect 1484 -7157 1517 -7086
rect 1550 -7129 1583 -7086
rect 1616 -7157 1649 -7086
rect 1682 -7129 1715 -7086
rect 1748 -7157 1781 -7086
rect 1814 -7129 1847 -7086
rect 1946 -7129 1979 -7086
rect 1880 -7157 1913 -7086
rect 1022 -7200 1055 -7157
rect 924 -7200 1022 -7157
rect 1022 -7200 1055 -7157
rect 1088 -7228 1121 -7157
rect 1154 -7200 1187 -7157
rect 1220 -7228 1253 -7157
rect 1286 -7200 1319 -7157
rect 1352 -7228 1385 -7157
rect 1418 -7200 1451 -7157
rect 1484 -7228 1517 -7157
rect 1550 -7200 1583 -7157
rect 1616 -7228 1649 -7157
rect 1682 -7200 1715 -7157
rect 1748 -7228 1781 -7157
rect 1814 -7200 1847 -7157
rect 1946 -7200 1979 -7157
rect 1880 -7228 1913 -7157
rect 1022 -7271 1055 -7228
rect 924 -7271 1022 -7228
rect 1022 -7271 1055 -7228
rect 1088 -7299 1121 -7228
rect 1154 -7271 1187 -7228
rect 1220 -7299 1253 -7228
rect 1286 -7271 1319 -7228
rect 1352 -7299 1385 -7228
rect 1418 -7271 1451 -7228
rect 1484 -7299 1517 -7228
rect 1550 -7271 1583 -7228
rect 1616 -7299 1649 -7228
rect 1682 -7271 1715 -7228
rect 1748 -7299 1781 -7228
rect 1814 -7271 1847 -7228
rect 1946 -7271 1979 -7228
rect 1880 -7299 1913 -7228
rect 1022 -7342 1055 -7299
rect 924 -7342 1022 -7299
rect 1022 -7342 1055 -7299
rect 1088 -7370 1121 -7299
rect 1154 -7342 1187 -7299
rect 1220 -7370 1253 -7299
rect 1286 -7342 1319 -7299
rect 1352 -7370 1385 -7299
rect 1418 -7342 1451 -7299
rect 1484 -7370 1517 -7299
rect 1550 -7342 1583 -7299
rect 1616 -7370 1649 -7299
rect 1682 -7342 1715 -7299
rect 1748 -7370 1781 -7299
rect 1814 -7342 1847 -7299
rect 1946 -7342 1979 -7299
rect 1880 -7370 1913 -7299
rect 1022 -7413 1055 -7370
rect 924 -7413 1022 -7370
rect 1022 -7413 1055 -7370
rect 1088 -7441 1121 -7370
rect 1154 -7413 1187 -7370
rect 1220 -7441 1253 -7370
rect 1286 -7413 1319 -7370
rect 1352 -7441 1385 -7370
rect 1418 -7413 1451 -7370
rect 1484 -7441 1517 -7370
rect 1550 -7413 1583 -7370
rect 1616 -7441 1649 -7370
rect 1682 -7413 1715 -7370
rect 1748 -7441 1781 -7370
rect 1814 -7413 1847 -7370
rect 1946 -7413 1979 -7370
rect 1880 -7441 1913 -7370
rect 1022 -7484 1055 -7441
rect 924 -7484 1022 -7441
rect 1022 -7484 1055 -7441
rect 1088 -7512 1121 -7441
rect 1154 -7484 1187 -7441
rect 1220 -7512 1253 -7441
rect 1286 -7484 1319 -7441
rect 1352 -7512 1385 -7441
rect 1418 -7484 1451 -7441
rect 1484 -7512 1517 -7441
rect 1550 -7484 1583 -7441
rect 1616 -7512 1649 -7441
rect 1682 -7484 1715 -7441
rect 1748 -7512 1781 -7441
rect 1814 -7484 1847 -7441
rect 1946 -7484 1979 -7441
rect 1880 -7512 1913 -7441
rect 1022 -7555 1055 -7512
rect 924 -7555 1022 -7512
rect 1022 -7555 1055 -7512
rect 1088 -7583 1121 -7512
rect 1154 -7555 1187 -7512
rect 1220 -7583 1253 -7512
rect 1286 -7555 1319 -7512
rect 1352 -7583 1385 -7512
rect 1418 -7555 1451 -7512
rect 1484 -7583 1517 -7512
rect 1550 -7555 1583 -7512
rect 1616 -7583 1649 -7512
rect 1682 -7555 1715 -7512
rect 1748 -7583 1781 -7512
rect 1814 -7555 1847 -7512
rect 1946 -7555 1979 -7512
rect 1880 -7583 1913 -7512
rect 1022 -7626 1055 -7583
rect 924 -7626 1022 -7583
rect 1022 -7626 1055 -7583
rect 1088 -7654 1121 -7583
rect 1154 -7626 1187 -7583
rect 1220 -7654 1253 -7583
rect 1286 -7626 1319 -7583
rect 1352 -7654 1385 -7583
rect 1418 -7626 1451 -7583
rect 1484 -7654 1517 -7583
rect 1550 -7626 1583 -7583
rect 1616 -7654 1649 -7583
rect 1682 -7626 1715 -7583
rect 1748 -7654 1781 -7583
rect 1814 -7626 1847 -7583
rect 1946 -7626 1979 -7583
rect 1880 -7654 1913 -7583
rect 1022 -7697 1055 -7654
rect 924 -7697 1022 -7654
rect 1022 -7697 1055 -7654
rect 1088 -7725 1121 -7654
rect 1154 -7697 1187 -7654
rect 1220 -7725 1253 -7654
rect 1286 -7697 1319 -7654
rect 1352 -7725 1385 -7654
rect 1418 -7697 1451 -7654
rect 1484 -7725 1517 -7654
rect 1550 -7697 1583 -7654
rect 1616 -7725 1649 -7654
rect 1682 -7697 1715 -7654
rect 1748 -7725 1781 -7654
rect 1814 -7697 1847 -7654
rect 1946 -7697 1979 -7654
rect 1880 -7725 1913 -7654
rect 1022 -7768 1055 -7725
rect 924 -7768 1022 -7725
rect 1022 -7768 1055 -7725
rect 1088 -7796 1121 -7725
rect 1154 -7768 1187 -7725
rect 1220 -7796 1253 -7725
rect 1286 -7768 1319 -7725
rect 1352 -7796 1385 -7725
rect 1418 -7768 1451 -7725
rect 1484 -7796 1517 -7725
rect 1550 -7768 1583 -7725
rect 1616 -7796 1649 -7725
rect 1682 -7768 1715 -7725
rect 1748 -7796 1781 -7725
rect 1814 -7768 1847 -7725
rect 1946 -7768 1979 -7725
rect 1880 -7796 1913 -7725
rect 1022 -7839 1055 -7796
rect 924 -7839 1022 -7796
rect 1022 -7839 1055 -7796
rect 1088 -7867 1121 -7796
rect 1154 -7839 1187 -7796
rect 1220 -7867 1253 -7796
rect 1286 -7839 1319 -7796
rect 1352 -7867 1385 -7796
rect 1418 -7839 1451 -7796
rect 1484 -7867 1517 -7796
rect 1550 -7839 1583 -7796
rect 1616 -7867 1649 -7796
rect 1682 -7839 1715 -7796
rect 1748 -7867 1781 -7796
rect 1814 -7839 1847 -7796
rect 1946 -7839 1979 -7796
rect 1880 -7867 1913 -7796
rect 1022 -7910 1055 -7867
rect 924 -7910 1022 -7867
rect 1022 -7910 1055 -7867
rect 1088 -7938 1121 -7867
rect 1154 -7910 1187 -7867
rect 1220 -7938 1253 -7867
rect 1286 -7910 1319 -7867
rect 1352 -7938 1385 -7867
rect 1418 -7910 1451 -7867
rect 1484 -7938 1517 -7867
rect 1550 -7910 1583 -7867
rect 1616 -7938 1649 -7867
rect 1682 -7910 1715 -7867
rect 1748 -7938 1781 -7867
rect 1814 -7910 1847 -7867
rect 1946 -7910 1979 -7867
rect 1880 -7938 1913 -7867
rect 1022 -7981 1055 -7938
rect 924 -7981 1022 -7938
rect 1022 -7981 1055 -7938
rect 1088 -8009 1121 -7938
rect 1154 -7981 1187 -7938
rect 1220 -8009 1253 -7938
rect 1286 -7981 1319 -7938
rect 1352 -8009 1385 -7938
rect 1418 -7981 1451 -7938
rect 1484 -8009 1517 -7938
rect 1550 -7981 1583 -7938
rect 1616 -8009 1649 -7938
rect 1682 -7981 1715 -7938
rect 1748 -8009 1781 -7938
rect 1814 -7981 1847 -7938
rect 1946 -7981 1979 -7938
rect 1880 -8009 1913 -7938
rect 1022 -8052 1055 -8009
rect 924 -8052 1022 -8009
rect 1022 -8052 1055 -8009
rect 1088 -8080 1121 -8009
rect 1154 -8052 1187 -8009
rect 1220 -8080 1253 -8009
rect 1286 -8052 1319 -8009
rect 1352 -8080 1385 -8009
rect 1418 -8052 1451 -8009
rect 1484 -8080 1517 -8009
rect 1550 -8052 1583 -8009
rect 1616 -8080 1649 -8009
rect 1682 -8052 1715 -8009
rect 1748 -8080 1781 -8009
rect 1814 -8052 1847 -8009
rect 1946 -8052 1979 -8009
rect 1880 -8080 1913 -8009
rect 1022 -8123 1055 -8080
rect 924 -8123 1022 -8080
rect 1022 -8123 1055 -8080
rect 1088 -8151 1121 -8080
rect 1154 -8123 1187 -8080
rect 1220 -8151 1253 -8080
rect 1286 -8123 1319 -8080
rect 1352 -8151 1385 -8080
rect 1418 -8123 1451 -8080
rect 1484 -8151 1517 -8080
rect 1550 -8123 1583 -8080
rect 1616 -8151 1649 -8080
rect 1682 -8123 1715 -8080
rect 1748 -8151 1781 -8080
rect 1814 -8123 1847 -8080
rect 1946 -8123 1979 -8080
rect 1880 -8151 1913 -8080
rect 1022 -8194 1055 -8151
rect 924 -8194 1022 -8151
rect 1022 -8194 1055 -8151
rect 1088 -8222 1121 -8151
rect 1154 -8194 1187 -8151
rect 1220 -8222 1253 -8151
rect 1286 -8194 1319 -8151
rect 1352 -8222 1385 -8151
rect 1418 -8194 1451 -8151
rect 1484 -8222 1517 -8151
rect 1550 -8194 1583 -8151
rect 1616 -8222 1649 -8151
rect 1682 -8194 1715 -8151
rect 1748 -8222 1781 -8151
rect 1814 -8194 1847 -8151
rect 1946 -8194 1979 -8151
rect 1880 -8222 1913 -8151
rect 1022 -8265 1055 -8222
rect 924 -8265 1022 -8222
rect 1022 -8265 1055 -8222
rect 1088 -8293 1121 -8222
rect 1154 -8265 1187 -8222
rect 1220 -8293 1253 -8222
rect 1286 -8265 1319 -8222
rect 1352 -8293 1385 -8222
rect 1418 -8265 1451 -8222
rect 1484 -8293 1517 -8222
rect 1550 -8265 1583 -8222
rect 1616 -8293 1649 -8222
rect 1682 -8265 1715 -8222
rect 1748 -8293 1781 -8222
rect 1814 -8265 1847 -8222
rect 1946 -8265 1979 -8222
rect 1880 -8293 1913 -8222
rect 1022 -8336 1055 -8293
rect 924 -8336 1022 -8293
rect 1022 -8336 1055 -8293
rect 1088 -8364 1121 -8293
rect 1154 -8336 1187 -8293
rect 1220 -8364 1253 -8293
rect 1286 -8336 1319 -8293
rect 1352 -8364 1385 -8293
rect 1418 -8336 1451 -8293
rect 1484 -8364 1517 -8293
rect 1550 -8336 1583 -8293
rect 1616 -8364 1649 -8293
rect 1682 -8336 1715 -8293
rect 1748 -8364 1781 -8293
rect 1814 -8336 1847 -8293
rect 1946 -8336 1979 -8293
rect 1880 -8364 1913 -8293
rect 1022 -8407 1055 -8364
rect 924 -8407 1022 -8364
rect 1022 -8407 1055 -8364
rect 1088 -8435 1121 -8364
rect 1154 -8407 1187 -8364
rect 1220 -8435 1253 -8364
rect 1286 -8407 1319 -8364
rect 1352 -8435 1385 -8364
rect 1418 -8407 1451 -8364
rect 1484 -8435 1517 -8364
rect 1550 -8407 1583 -8364
rect 1616 -8435 1649 -8364
rect 1682 -8407 1715 -8364
rect 1748 -8435 1781 -8364
rect 1814 -8407 1847 -8364
rect 1946 -8407 1979 -8364
rect 1880 -8435 1913 -8364
rect 1022 -8478 1055 -8435
rect 924 -8478 1022 -8435
rect 1022 -8478 1055 -8435
rect 1088 -8506 1121 -8435
rect 1154 -8478 1187 -8435
rect 1220 -8506 1253 -8435
rect 1286 -8478 1319 -8435
rect 1352 -8506 1385 -8435
rect 1418 -8478 1451 -8435
rect 1484 -8506 1517 -8435
rect 1550 -8478 1583 -8435
rect 1616 -8506 1649 -8435
rect 1682 -8478 1715 -8435
rect 1748 -8506 1781 -8435
rect 1814 -8478 1847 -8435
rect 1946 -8478 1979 -8435
rect 1880 -8506 1913 -8435
rect 1022 -8549 1055 -8506
rect 924 -8549 1022 -8506
rect 1022 -8549 1055 -8506
rect 1088 -8577 1121 -8506
rect 1154 -8549 1187 -8506
rect 1220 -8577 1253 -8506
rect 1286 -8549 1319 -8506
rect 1352 -8577 1385 -8506
rect 1418 -8549 1451 -8506
rect 1484 -8577 1517 -8506
rect 1550 -8549 1583 -8506
rect 1616 -8577 1649 -8506
rect 1682 -8549 1715 -8506
rect 1748 -8577 1781 -8506
rect 1814 -8549 1847 -8506
rect 1946 -8549 1979 -8506
rect 1880 -8577 1913 -8506
rect 1022 -8620 1055 -8577
rect 924 -8620 1022 -8577
rect 1022 -8620 1055 -8577
rect 1088 -8648 1121 -8577
rect 1154 -8620 1187 -8577
rect 1220 -8648 1253 -8577
rect 1286 -8620 1319 -8577
rect 1352 -8648 1385 -8577
rect 1418 -8620 1451 -8577
rect 1484 -8648 1517 -8577
rect 1550 -8620 1583 -8577
rect 1616 -8648 1649 -8577
rect 1682 -8620 1715 -8577
rect 1748 -8648 1781 -8577
rect 1814 -8620 1847 -8577
rect 1946 -8620 1979 -8577
rect 1880 -8648 1913 -8577
rect 1022 -8691 1055 -8648
rect 924 -8691 1022 -8648
rect 1022 -8691 1055 -8648
rect 1088 -8719 1121 -8648
rect 1154 -8691 1187 -8648
rect 1220 -8719 1253 -8648
rect 1286 -8691 1319 -8648
rect 1352 -8719 1385 -8648
rect 1418 -8691 1451 -8648
rect 1484 -8719 1517 -8648
rect 1550 -8691 1583 -8648
rect 1616 -8719 1649 -8648
rect 1682 -8691 1715 -8648
rect 1748 -8719 1781 -8648
rect 1814 -8691 1847 -8648
rect 1946 -8691 1979 -8648
rect 1880 -8719 1913 -8648
rect 1022 -8762 1055 -8719
rect 924 -8762 1022 -8719
rect 1022 -8762 1055 -8719
rect 1088 -8790 1121 -8719
rect 1154 -8762 1187 -8719
rect 1220 -8790 1253 -8719
rect 1286 -8762 1319 -8719
rect 1352 -8790 1385 -8719
rect 1418 -8762 1451 -8719
rect 1484 -8790 1517 -8719
rect 1550 -8762 1583 -8719
rect 1616 -8790 1649 -8719
rect 1682 -8762 1715 -8719
rect 1748 -8790 1781 -8719
rect 1814 -8762 1847 -8719
rect 1946 -8762 1979 -8719
rect 1880 -8790 1913 -8719
rect 1022 -8833 1055 -8790
rect 924 -8833 1022 -8790
rect 1022 -8833 1055 -8790
rect 1088 -8861 1121 -8790
rect 1154 -8833 1187 -8790
rect 1220 -8861 1253 -8790
rect 1286 -8833 1319 -8790
rect 1352 -8861 1385 -8790
rect 1418 -8833 1451 -8790
rect 1484 -8861 1517 -8790
rect 1550 -8833 1583 -8790
rect 1616 -8861 1649 -8790
rect 1682 -8833 1715 -8790
rect 1748 -8861 1781 -8790
rect 1814 -8833 1847 -8790
rect 1946 -8833 1979 -8790
rect 1880 -8861 1913 -8790
rect 1022 -8904 1055 -8861
rect 924 -8904 1022 -8861
rect 1022 -8904 1055 -8861
rect 1088 -8932 1121 -8861
rect 1154 -8904 1187 -8861
rect 1220 -8932 1253 -8861
rect 1286 -8904 1319 -8861
rect 1352 -8932 1385 -8861
rect 1418 -8904 1451 -8861
rect 1484 -8932 1517 -8861
rect 1550 -8904 1583 -8861
rect 1616 -8932 1649 -8861
rect 1682 -8904 1715 -8861
rect 1748 -8932 1781 -8861
rect 1814 -8904 1847 -8861
rect 1946 -8904 1979 -8861
rect 1880 -8932 1913 -8861
rect 1022 -8975 1055 -8932
rect 924 -8975 1022 -8932
rect 1022 -8975 1055 -8932
rect 1088 -9003 1121 -8932
rect 1154 -8975 1187 -8932
rect 1220 -9003 1253 -8932
rect 1286 -8975 1319 -8932
rect 1352 -9003 1385 -8932
rect 1418 -8975 1451 -8932
rect 1484 -9003 1517 -8932
rect 1550 -8975 1583 -8932
rect 1616 -9003 1649 -8932
rect 1682 -8975 1715 -8932
rect 1748 -9003 1781 -8932
rect 1814 -8975 1847 -8932
rect 1946 -8975 1979 -8932
rect 1880 -9003 1913 -8932
rect 1022 -9046 1055 -9003
rect 924 -9046 1022 -9003
rect 1022 -9046 1055 -9003
rect 1088 -9074 1121 -9003
rect 1154 -9046 1187 -9003
rect 1220 -9074 1253 -9003
rect 1286 -9046 1319 -9003
rect 1352 -9074 1385 -9003
rect 1418 -9046 1451 -9003
rect 1484 -9074 1517 -9003
rect 1550 -9046 1583 -9003
rect 1616 -9074 1649 -9003
rect 1682 -9046 1715 -9003
rect 1748 -9074 1781 -9003
rect 1814 -9046 1847 -9003
rect 1946 -9046 1979 -9003
rect 1880 -9074 1913 -9003
rect 1022 -9117 1055 -9074
rect 924 -9117 1022 -9074
rect 1022 -9117 1055 -9074
rect 1088 -9145 1121 -9074
rect 1154 -9117 1187 -9074
rect 1220 -9145 1253 -9074
rect 1286 -9117 1319 -9074
rect 1352 -9145 1385 -9074
rect 1418 -9117 1451 -9074
rect 1484 -9145 1517 -9074
rect 1550 -9117 1583 -9074
rect 1616 -9145 1649 -9074
rect 1682 -9117 1715 -9074
rect 1748 -9145 1781 -9074
rect 1814 -9117 1847 -9074
rect 1946 -9117 1979 -9074
rect 1880 -9145 1913 -9074
rect -101 17 1946 65
rect -101 252 1946 300
rect -101 -9145 -53 17
rect 1022 -9193 1979 -9145
rect 1979 -9193 2059 -9145
rect 2019 -9145 2059 300
rect 1946 252 2019 300
rect 56 65 89 125
rect 0 82 33 125
rect 0 82 33 192
rect 56 142 89 175
rect 0 192 33 235
rect 56 192 89 252
rect 188 65 221 125
rect 132 82 165 125
rect 132 82 165 192
rect 188 142 221 175
rect 132 192 165 235
rect 188 192 221 252
rect 320 65 353 125
rect 264 82 297 125
rect 264 82 297 192
rect 320 142 353 175
rect 264 192 297 235
rect 320 192 353 252
rect 452 65 485 125
rect 396 82 429 125
rect 396 82 429 192
rect 452 142 485 175
rect 396 192 429 235
rect 452 192 485 252
rect 584 65 617 125
rect 528 82 561 125
rect 528 82 561 192
rect 584 142 617 175
rect 528 192 561 235
rect 584 192 617 252
rect 716 65 749 125
rect 660 82 693 125
rect 660 82 693 192
rect 716 142 749 175
rect 660 192 693 235
rect 716 192 749 252
rect 848 65 881 125
rect 792 82 825 125
rect 792 82 825 192
rect 848 142 881 175
rect 792 192 825 235
rect 848 192 881 252
rect 1065 65 1098 125
rect 1121 82 1154 125
rect 1121 82 1154 192
rect 1065 142 1098 175
rect 1121 192 1154 235
rect 1065 192 1098 252
rect 1197 65 1230 125
rect 1253 82 1286 125
rect 1253 82 1286 192
rect 1197 142 1230 175
rect 1253 192 1286 235
rect 1197 192 1230 252
rect 1329 65 1362 125
rect 1385 82 1418 125
rect 1385 82 1418 192
rect 1329 142 1362 175
rect 1385 192 1418 235
rect 1329 192 1362 252
rect 1461 65 1494 125
rect 1517 82 1550 125
rect 1517 82 1550 192
rect 1461 142 1494 175
rect 1517 192 1550 235
rect 1461 192 1494 252
rect 1593 65 1626 125
rect 1649 82 1682 125
rect 1649 82 1682 192
rect 1593 142 1626 175
rect 1649 192 1682 235
rect 1593 192 1626 252
rect 1725 65 1758 125
rect 1781 82 1814 125
rect 1781 82 1814 192
rect 1725 142 1758 175
rect 1781 192 1814 235
rect 1725 192 1758 252
rect 1857 65 1890 125
rect 1913 82 1946 125
rect 1913 82 1946 192
rect 1857 142 1890 175
rect 1913 192 1946 235
rect 1857 192 1890 252
<< nwell >>
rect -119 -9147 942 143
rect 942 7 1948 143
<< viali >>
rect 8 -25 25 -8
rect 74 -25 91 -8
rect 140 -25 157 -8
rect 206 -25 223 -8
rect 272 -25 289 -8
rect 338 -25 355 -8
rect 404 -25 421 -8
rect 470 -25 487 -8
rect 536 -25 553 -8
rect 602 -25 619 -8
rect 668 -25 685 -8
rect 734 -25 751 -8
rect 800 -25 817 -8
rect 866 -25 883 -8
rect 1063 -25 1080 -8
rect 1129 -25 1146 -8
rect 1195 -25 1212 -8
rect 1261 -25 1278 -8
rect 1327 -25 1344 -8
rect 1393 -25 1410 -8
rect 1459 -25 1476 -8
rect 1525 -25 1542 -8
rect 1591 -25 1608 -8
rect 1657 -25 1674 -8
rect 1723 -25 1740 -8
rect 1789 -25 1806 -8
rect 1855 -25 1872 -8
rect 1921 -25 1938 -8
rect 1030 -92 1047 -65
rect 1030 -92 1047 -65
rect 1162 -92 1179 -65
rect 1294 -92 1311 -65
rect 1426 -92 1443 -65
rect 1558 -92 1575 -65
rect 1690 -92 1707 -65
rect 1822 -92 1839 -65
rect 1030 -163 1047 -136
rect 1030 -163 1047 -136
rect 1162 -163 1179 -136
rect 1294 -163 1311 -136
rect 1426 -163 1443 -136
rect 1558 -163 1575 -136
rect 1690 -163 1707 -136
rect 1822 -163 1839 -136
rect 1030 -234 1047 -207
rect 1030 -234 1047 -207
rect 1162 -234 1179 -207
rect 1294 -234 1311 -207
rect 1426 -234 1443 -207
rect 1558 -234 1575 -207
rect 1690 -234 1707 -207
rect 1822 -234 1839 -207
rect 1030 -305 1047 -278
rect 1030 -305 1047 -278
rect 1162 -305 1179 -278
rect 1294 -305 1311 -278
rect 1426 -305 1443 -278
rect 1558 -305 1575 -278
rect 1690 -305 1707 -278
rect 1822 -305 1839 -278
rect 1030 -376 1047 -349
rect 1030 -376 1047 -349
rect 1162 -376 1179 -349
rect 1294 -376 1311 -349
rect 1426 -376 1443 -349
rect 1558 -376 1575 -349
rect 1690 -376 1707 -349
rect 1822 -376 1839 -349
rect 1030 -447 1047 -420
rect 1030 -447 1047 -420
rect 1162 -447 1179 -420
rect 1294 -447 1311 -420
rect 1426 -447 1443 -420
rect 1558 -447 1575 -420
rect 1690 -447 1707 -420
rect 1822 -447 1839 -420
rect 1030 -518 1047 -491
rect 1030 -518 1047 -491
rect 1162 -518 1179 -491
rect 1294 -518 1311 -491
rect 1426 -518 1443 -491
rect 1558 -518 1575 -491
rect 1690 -518 1707 -491
rect 1822 -518 1839 -491
rect 1030 -589 1047 -562
rect 1030 -589 1047 -562
rect 1162 -589 1179 -562
rect 1294 -589 1311 -562
rect 1426 -589 1443 -562
rect 1558 -589 1575 -562
rect 1690 -589 1707 -562
rect 1822 -589 1839 -562
rect 1030 -660 1047 -633
rect 1030 -660 1047 -633
rect 1162 -660 1179 -633
rect 1294 -660 1311 -633
rect 1426 -660 1443 -633
rect 1558 -660 1575 -633
rect 1690 -660 1707 -633
rect 1822 -660 1839 -633
rect 1030 -731 1047 -704
rect 1030 -731 1047 -704
rect 1162 -731 1179 -704
rect 1294 -731 1311 -704
rect 1426 -731 1443 -704
rect 1558 -731 1575 -704
rect 1690 -731 1707 -704
rect 1822 -731 1839 -704
rect 1030 -802 1047 -775
rect 1030 -802 1047 -775
rect 1162 -802 1179 -775
rect 1294 -802 1311 -775
rect 1426 -802 1443 -775
rect 1558 -802 1575 -775
rect 1690 -802 1707 -775
rect 1822 -802 1839 -775
rect 1030 -873 1047 -846
rect 1030 -873 1047 -846
rect 1162 -873 1179 -846
rect 1294 -873 1311 -846
rect 1426 -873 1443 -846
rect 1558 -873 1575 -846
rect 1690 -873 1707 -846
rect 1822 -873 1839 -846
rect 1030 -944 1047 -917
rect 1030 -944 1047 -917
rect 1162 -944 1179 -917
rect 1294 -944 1311 -917
rect 1426 -944 1443 -917
rect 1558 -944 1575 -917
rect 1690 -944 1707 -917
rect 1822 -944 1839 -917
rect 1030 -1015 1047 -988
rect 1030 -1015 1047 -988
rect 1162 -1015 1179 -988
rect 1294 -1015 1311 -988
rect 1426 -1015 1443 -988
rect 1558 -1015 1575 -988
rect 1690 -1015 1707 -988
rect 1822 -1015 1839 -988
rect 1030 -1086 1047 -1059
rect 1030 -1086 1047 -1059
rect 1162 -1086 1179 -1059
rect 1294 -1086 1311 -1059
rect 1426 -1086 1443 -1059
rect 1558 -1086 1575 -1059
rect 1690 -1086 1707 -1059
rect 1822 -1086 1839 -1059
rect 1030 -1157 1047 -1130
rect 1030 -1157 1047 -1130
rect 1162 -1157 1179 -1130
rect 1294 -1157 1311 -1130
rect 1426 -1157 1443 -1130
rect 1558 -1157 1575 -1130
rect 1690 -1157 1707 -1130
rect 1822 -1157 1839 -1130
rect 1030 -1228 1047 -1201
rect 1030 -1228 1047 -1201
rect 1162 -1228 1179 -1201
rect 1294 -1228 1311 -1201
rect 1426 -1228 1443 -1201
rect 1558 -1228 1575 -1201
rect 1690 -1228 1707 -1201
rect 1822 -1228 1839 -1201
rect 1030 -1299 1047 -1272
rect 1030 -1299 1047 -1272
rect 1162 -1299 1179 -1272
rect 1294 -1299 1311 -1272
rect 1426 -1299 1443 -1272
rect 1558 -1299 1575 -1272
rect 1690 -1299 1707 -1272
rect 1822 -1299 1839 -1272
rect 1030 -1370 1047 -1343
rect 1030 -1370 1047 -1343
rect 1162 -1370 1179 -1343
rect 1294 -1370 1311 -1343
rect 1426 -1370 1443 -1343
rect 1558 -1370 1575 -1343
rect 1690 -1370 1707 -1343
rect 1822 -1370 1839 -1343
rect 1030 -1441 1047 -1414
rect 1030 -1441 1047 -1414
rect 1162 -1441 1179 -1414
rect 1294 -1441 1311 -1414
rect 1426 -1441 1443 -1414
rect 1558 -1441 1575 -1414
rect 1690 -1441 1707 -1414
rect 1822 -1441 1839 -1414
rect 1030 -1512 1047 -1485
rect 1030 -1512 1047 -1485
rect 1162 -1512 1179 -1485
rect 1294 -1512 1311 -1485
rect 1426 -1512 1443 -1485
rect 1558 -1512 1575 -1485
rect 1690 -1512 1707 -1485
rect 1822 -1512 1839 -1485
rect 1030 -1583 1047 -1556
rect 1030 -1583 1047 -1556
rect 1162 -1583 1179 -1556
rect 1294 -1583 1311 -1556
rect 1426 -1583 1443 -1556
rect 1558 -1583 1575 -1556
rect 1690 -1583 1707 -1556
rect 1822 -1583 1839 -1556
rect 1030 -1654 1047 -1627
rect 1030 -1654 1047 -1627
rect 1162 -1654 1179 -1627
rect 1294 -1654 1311 -1627
rect 1426 -1654 1443 -1627
rect 1558 -1654 1575 -1627
rect 1690 -1654 1707 -1627
rect 1822 -1654 1839 -1627
rect 1030 -1725 1047 -1698
rect 1030 -1725 1047 -1698
rect 1162 -1725 1179 -1698
rect 1294 -1725 1311 -1698
rect 1426 -1725 1443 -1698
rect 1558 -1725 1575 -1698
rect 1690 -1725 1707 -1698
rect 1822 -1725 1839 -1698
rect 1030 -1796 1047 -1769
rect 1030 -1796 1047 -1769
rect 1162 -1796 1179 -1769
rect 1294 -1796 1311 -1769
rect 1426 -1796 1443 -1769
rect 1558 -1796 1575 -1769
rect 1690 -1796 1707 -1769
rect 1822 -1796 1839 -1769
rect 1030 -1867 1047 -1840
rect 1030 -1867 1047 -1840
rect 1162 -1867 1179 -1840
rect 1294 -1867 1311 -1840
rect 1426 -1867 1443 -1840
rect 1558 -1867 1575 -1840
rect 1690 -1867 1707 -1840
rect 1822 -1867 1839 -1840
rect 1030 -1938 1047 -1911
rect 1030 -1938 1047 -1911
rect 1162 -1938 1179 -1911
rect 1294 -1938 1311 -1911
rect 1426 -1938 1443 -1911
rect 1558 -1938 1575 -1911
rect 1690 -1938 1707 -1911
rect 1822 -1938 1839 -1911
rect 1030 -2009 1047 -1982
rect 1030 -2009 1047 -1982
rect 1162 -2009 1179 -1982
rect 1294 -2009 1311 -1982
rect 1426 -2009 1443 -1982
rect 1558 -2009 1575 -1982
rect 1690 -2009 1707 -1982
rect 1822 -2009 1839 -1982
rect 1030 -2080 1047 -2053
rect 1030 -2080 1047 -2053
rect 1162 -2080 1179 -2053
rect 1294 -2080 1311 -2053
rect 1426 -2080 1443 -2053
rect 1558 -2080 1575 -2053
rect 1690 -2080 1707 -2053
rect 1822 -2080 1839 -2053
rect 1030 -2151 1047 -2124
rect 1030 -2151 1047 -2124
rect 1162 -2151 1179 -2124
rect 1294 -2151 1311 -2124
rect 1426 -2151 1443 -2124
rect 1558 -2151 1575 -2124
rect 1690 -2151 1707 -2124
rect 1822 -2151 1839 -2124
rect 1030 -2222 1047 -2195
rect 1030 -2222 1047 -2195
rect 1162 -2222 1179 -2195
rect 1294 -2222 1311 -2195
rect 1426 -2222 1443 -2195
rect 1558 -2222 1575 -2195
rect 1690 -2222 1707 -2195
rect 1822 -2222 1839 -2195
rect 1030 -2293 1047 -2266
rect 1030 -2293 1047 -2266
rect 1162 -2293 1179 -2266
rect 1294 -2293 1311 -2266
rect 1426 -2293 1443 -2266
rect 1558 -2293 1575 -2266
rect 1690 -2293 1707 -2266
rect 1822 -2293 1839 -2266
rect 1030 -2364 1047 -2337
rect 1030 -2364 1047 -2337
rect 1162 -2364 1179 -2337
rect 1294 -2364 1311 -2337
rect 1426 -2364 1443 -2337
rect 1558 -2364 1575 -2337
rect 1690 -2364 1707 -2337
rect 1822 -2364 1839 -2337
rect 1030 -2435 1047 -2408
rect 1030 -2435 1047 -2408
rect 1162 -2435 1179 -2408
rect 1294 -2435 1311 -2408
rect 1426 -2435 1443 -2408
rect 1558 -2435 1575 -2408
rect 1690 -2435 1707 -2408
rect 1822 -2435 1839 -2408
rect 1030 -2506 1047 -2479
rect 1030 -2506 1047 -2479
rect 1162 -2506 1179 -2479
rect 1294 -2506 1311 -2479
rect 1426 -2506 1443 -2479
rect 1558 -2506 1575 -2479
rect 1690 -2506 1707 -2479
rect 1822 -2506 1839 -2479
rect 1030 -2577 1047 -2550
rect 1030 -2577 1047 -2550
rect 1162 -2577 1179 -2550
rect 1294 -2577 1311 -2550
rect 1426 -2577 1443 -2550
rect 1558 -2577 1575 -2550
rect 1690 -2577 1707 -2550
rect 1822 -2577 1839 -2550
rect 1030 -2648 1047 -2621
rect 1030 -2648 1047 -2621
rect 1162 -2648 1179 -2621
rect 1294 -2648 1311 -2621
rect 1426 -2648 1443 -2621
rect 1558 -2648 1575 -2621
rect 1690 -2648 1707 -2621
rect 1822 -2648 1839 -2621
rect 1030 -2719 1047 -2692
rect 1030 -2719 1047 -2692
rect 1162 -2719 1179 -2692
rect 1294 -2719 1311 -2692
rect 1426 -2719 1443 -2692
rect 1558 -2719 1575 -2692
rect 1690 -2719 1707 -2692
rect 1822 -2719 1839 -2692
rect 1030 -2790 1047 -2763
rect 1030 -2790 1047 -2763
rect 1162 -2790 1179 -2763
rect 1294 -2790 1311 -2763
rect 1426 -2790 1443 -2763
rect 1558 -2790 1575 -2763
rect 1690 -2790 1707 -2763
rect 1822 -2790 1839 -2763
rect 1030 -2861 1047 -2834
rect 1030 -2861 1047 -2834
rect 1162 -2861 1179 -2834
rect 1294 -2861 1311 -2834
rect 1426 -2861 1443 -2834
rect 1558 -2861 1575 -2834
rect 1690 -2861 1707 -2834
rect 1822 -2861 1839 -2834
rect 1030 -2932 1047 -2905
rect 1030 -2932 1047 -2905
rect 1162 -2932 1179 -2905
rect 1294 -2932 1311 -2905
rect 1426 -2932 1443 -2905
rect 1558 -2932 1575 -2905
rect 1690 -2932 1707 -2905
rect 1822 -2932 1839 -2905
rect 1030 -3003 1047 -2976
rect 1030 -3003 1047 -2976
rect 1162 -3003 1179 -2976
rect 1294 -3003 1311 -2976
rect 1426 -3003 1443 -2976
rect 1558 -3003 1575 -2976
rect 1690 -3003 1707 -2976
rect 1822 -3003 1839 -2976
rect 1030 -3074 1047 -3047
rect 1030 -3074 1047 -3047
rect 1162 -3074 1179 -3047
rect 1294 -3074 1311 -3047
rect 1426 -3074 1443 -3047
rect 1558 -3074 1575 -3047
rect 1690 -3074 1707 -3047
rect 1822 -3074 1839 -3047
rect 1030 -3145 1047 -3118
rect 1030 -3145 1047 -3118
rect 1162 -3145 1179 -3118
rect 1294 -3145 1311 -3118
rect 1426 -3145 1443 -3118
rect 1558 -3145 1575 -3118
rect 1690 -3145 1707 -3118
rect 1822 -3145 1839 -3118
rect 1030 -3216 1047 -3189
rect 1030 -3216 1047 -3189
rect 1162 -3216 1179 -3189
rect 1294 -3216 1311 -3189
rect 1426 -3216 1443 -3189
rect 1558 -3216 1575 -3189
rect 1690 -3216 1707 -3189
rect 1822 -3216 1839 -3189
rect 1030 -3287 1047 -3260
rect 1030 -3287 1047 -3260
rect 1162 -3287 1179 -3260
rect 1294 -3287 1311 -3260
rect 1426 -3287 1443 -3260
rect 1558 -3287 1575 -3260
rect 1690 -3287 1707 -3260
rect 1822 -3287 1839 -3260
rect 1030 -3358 1047 -3331
rect 1030 -3358 1047 -3331
rect 1162 -3358 1179 -3331
rect 1294 -3358 1311 -3331
rect 1426 -3358 1443 -3331
rect 1558 -3358 1575 -3331
rect 1690 -3358 1707 -3331
rect 1822 -3358 1839 -3331
rect 1030 -3429 1047 -3402
rect 1030 -3429 1047 -3402
rect 1162 -3429 1179 -3402
rect 1294 -3429 1311 -3402
rect 1426 -3429 1443 -3402
rect 1558 -3429 1575 -3402
rect 1690 -3429 1707 -3402
rect 1822 -3429 1839 -3402
rect 1030 -3500 1047 -3473
rect 1030 -3500 1047 -3473
rect 1162 -3500 1179 -3473
rect 1294 -3500 1311 -3473
rect 1426 -3500 1443 -3473
rect 1558 -3500 1575 -3473
rect 1690 -3500 1707 -3473
rect 1822 -3500 1839 -3473
rect 1030 -3571 1047 -3544
rect 1030 -3571 1047 -3544
rect 1162 -3571 1179 -3544
rect 1294 -3571 1311 -3544
rect 1426 -3571 1443 -3544
rect 1558 -3571 1575 -3544
rect 1690 -3571 1707 -3544
rect 1822 -3571 1839 -3544
rect 1030 -3642 1047 -3615
rect 1030 -3642 1047 -3615
rect 1162 -3642 1179 -3615
rect 1294 -3642 1311 -3615
rect 1426 -3642 1443 -3615
rect 1558 -3642 1575 -3615
rect 1690 -3642 1707 -3615
rect 1822 -3642 1839 -3615
rect 1030 -3713 1047 -3686
rect 1030 -3713 1047 -3686
rect 1162 -3713 1179 -3686
rect 1294 -3713 1311 -3686
rect 1426 -3713 1443 -3686
rect 1558 -3713 1575 -3686
rect 1690 -3713 1707 -3686
rect 1822 -3713 1839 -3686
rect 1030 -3784 1047 -3757
rect 1030 -3784 1047 -3757
rect 1162 -3784 1179 -3757
rect 1294 -3784 1311 -3757
rect 1426 -3784 1443 -3757
rect 1558 -3784 1575 -3757
rect 1690 -3784 1707 -3757
rect 1822 -3784 1839 -3757
rect 1030 -3855 1047 -3828
rect 1030 -3855 1047 -3828
rect 1162 -3855 1179 -3828
rect 1294 -3855 1311 -3828
rect 1426 -3855 1443 -3828
rect 1558 -3855 1575 -3828
rect 1690 -3855 1707 -3828
rect 1822 -3855 1839 -3828
rect 1030 -3926 1047 -3899
rect 1030 -3926 1047 -3899
rect 1162 -3926 1179 -3899
rect 1294 -3926 1311 -3899
rect 1426 -3926 1443 -3899
rect 1558 -3926 1575 -3899
rect 1690 -3926 1707 -3899
rect 1822 -3926 1839 -3899
rect 1030 -3997 1047 -3970
rect 1030 -3997 1047 -3970
rect 1162 -3997 1179 -3970
rect 1294 -3997 1311 -3970
rect 1426 -3997 1443 -3970
rect 1558 -3997 1575 -3970
rect 1690 -3997 1707 -3970
rect 1822 -3997 1839 -3970
rect 1030 -4068 1047 -4041
rect 1030 -4068 1047 -4041
rect 1162 -4068 1179 -4041
rect 1294 -4068 1311 -4041
rect 1426 -4068 1443 -4041
rect 1558 -4068 1575 -4041
rect 1690 -4068 1707 -4041
rect 1822 -4068 1839 -4041
rect 1030 -4139 1047 -4112
rect 1030 -4139 1047 -4112
rect 1162 -4139 1179 -4112
rect 1294 -4139 1311 -4112
rect 1426 -4139 1443 -4112
rect 1558 -4139 1575 -4112
rect 1690 -4139 1707 -4112
rect 1822 -4139 1839 -4112
rect 1030 -4210 1047 -4183
rect 1030 -4210 1047 -4183
rect 1162 -4210 1179 -4183
rect 1294 -4210 1311 -4183
rect 1426 -4210 1443 -4183
rect 1558 -4210 1575 -4183
rect 1690 -4210 1707 -4183
rect 1822 -4210 1839 -4183
rect 1030 -4281 1047 -4254
rect 1030 -4281 1047 -4254
rect 1162 -4281 1179 -4254
rect 1294 -4281 1311 -4254
rect 1426 -4281 1443 -4254
rect 1558 -4281 1575 -4254
rect 1690 -4281 1707 -4254
rect 1822 -4281 1839 -4254
rect 1030 -4352 1047 -4325
rect 1030 -4352 1047 -4325
rect 1162 -4352 1179 -4325
rect 1294 -4352 1311 -4325
rect 1426 -4352 1443 -4325
rect 1558 -4352 1575 -4325
rect 1690 -4352 1707 -4325
rect 1822 -4352 1839 -4325
rect 1030 -4423 1047 -4396
rect 1030 -4423 1047 -4396
rect 1162 -4423 1179 -4396
rect 1294 -4423 1311 -4396
rect 1426 -4423 1443 -4396
rect 1558 -4423 1575 -4396
rect 1690 -4423 1707 -4396
rect 1822 -4423 1839 -4396
rect 1030 -4494 1047 -4467
rect 1030 -4494 1047 -4467
rect 1162 -4494 1179 -4467
rect 1294 -4494 1311 -4467
rect 1426 -4494 1443 -4467
rect 1558 -4494 1575 -4467
rect 1690 -4494 1707 -4467
rect 1822 -4494 1839 -4467
rect 1030 -4565 1047 -4538
rect 1030 -4565 1047 -4538
rect 1162 -4565 1179 -4538
rect 1294 -4565 1311 -4538
rect 1426 -4565 1443 -4538
rect 1558 -4565 1575 -4538
rect 1690 -4565 1707 -4538
rect 1822 -4565 1839 -4538
rect 1030 -4636 1047 -4609
rect 1030 -4636 1047 -4609
rect 1162 -4636 1179 -4609
rect 1294 -4636 1311 -4609
rect 1426 -4636 1443 -4609
rect 1558 -4636 1575 -4609
rect 1690 -4636 1707 -4609
rect 1822 -4636 1839 -4609
rect 1954 -4636 1971 -4609
rect 1030 -4707 1047 -4680
rect 1030 -4707 1047 -4680
rect 1162 -4707 1179 -4680
rect 1294 -4707 1311 -4680
rect 1426 -4707 1443 -4680
rect 1558 -4707 1575 -4680
rect 1690 -4707 1707 -4680
rect 1822 -4707 1839 -4680
rect 1954 -4707 1971 -4680
rect 1030 -4778 1047 -4751
rect 1030 -4778 1047 -4751
rect 1162 -4778 1179 -4751
rect 1294 -4778 1311 -4751
rect 1426 -4778 1443 -4751
rect 1558 -4778 1575 -4751
rect 1690 -4778 1707 -4751
rect 1822 -4778 1839 -4751
rect 1954 -4778 1971 -4751
rect 1030 -4849 1047 -4822
rect 1030 -4849 1047 -4822
rect 1162 -4849 1179 -4822
rect 1294 -4849 1311 -4822
rect 1426 -4849 1443 -4822
rect 1558 -4849 1575 -4822
rect 1690 -4849 1707 -4822
rect 1822 -4849 1839 -4822
rect 1954 -4849 1971 -4822
rect 1030 -4920 1047 -4893
rect 1030 -4920 1047 -4893
rect 1162 -4920 1179 -4893
rect 1294 -4920 1311 -4893
rect 1426 -4920 1443 -4893
rect 1558 -4920 1575 -4893
rect 1690 -4920 1707 -4893
rect 1822 -4920 1839 -4893
rect 1954 -4920 1971 -4893
rect 1030 -4991 1047 -4964
rect 1030 -4991 1047 -4964
rect 1162 -4991 1179 -4964
rect 1294 -4991 1311 -4964
rect 1426 -4991 1443 -4964
rect 1558 -4991 1575 -4964
rect 1690 -4991 1707 -4964
rect 1822 -4991 1839 -4964
rect 1954 -4991 1971 -4964
rect 1030 -5062 1047 -5035
rect 1030 -5062 1047 -5035
rect 1162 -5062 1179 -5035
rect 1294 -5062 1311 -5035
rect 1426 -5062 1443 -5035
rect 1558 -5062 1575 -5035
rect 1690 -5062 1707 -5035
rect 1822 -5062 1839 -5035
rect 1954 -5062 1971 -5035
rect 1030 -5133 1047 -5106
rect 1030 -5133 1047 -5106
rect 1162 -5133 1179 -5106
rect 1294 -5133 1311 -5106
rect 1426 -5133 1443 -5106
rect 1558 -5133 1575 -5106
rect 1690 -5133 1707 -5106
rect 1822 -5133 1839 -5106
rect 1954 -5133 1971 -5106
rect 1030 -5204 1047 -5177
rect 1030 -5204 1047 -5177
rect 1162 -5204 1179 -5177
rect 1294 -5204 1311 -5177
rect 1426 -5204 1443 -5177
rect 1558 -5204 1575 -5177
rect 1690 -5204 1707 -5177
rect 1822 -5204 1839 -5177
rect 1954 -5204 1971 -5177
rect 1030 -5275 1047 -5248
rect 1030 -5275 1047 -5248
rect 1162 -5275 1179 -5248
rect 1294 -5275 1311 -5248
rect 1426 -5275 1443 -5248
rect 1558 -5275 1575 -5248
rect 1690 -5275 1707 -5248
rect 1822 -5275 1839 -5248
rect 1954 -5275 1971 -5248
rect 1030 -5346 1047 -5319
rect 1030 -5346 1047 -5319
rect 1162 -5346 1179 -5319
rect 1294 -5346 1311 -5319
rect 1426 -5346 1443 -5319
rect 1558 -5346 1575 -5319
rect 1690 -5346 1707 -5319
rect 1822 -5346 1839 -5319
rect 1954 -5346 1971 -5319
rect 1030 -5417 1047 -5390
rect 1030 -5417 1047 -5390
rect 1162 -5417 1179 -5390
rect 1294 -5417 1311 -5390
rect 1426 -5417 1443 -5390
rect 1558 -5417 1575 -5390
rect 1690 -5417 1707 -5390
rect 1822 -5417 1839 -5390
rect 1954 -5417 1971 -5390
rect 1030 -5488 1047 -5461
rect 1030 -5488 1047 -5461
rect 1162 -5488 1179 -5461
rect 1294 -5488 1311 -5461
rect 1426 -5488 1443 -5461
rect 1558 -5488 1575 -5461
rect 1690 -5488 1707 -5461
rect 1822 -5488 1839 -5461
rect 1954 -5488 1971 -5461
rect 1030 -5559 1047 -5532
rect 1030 -5559 1047 -5532
rect 1162 -5559 1179 -5532
rect 1294 -5559 1311 -5532
rect 1426 -5559 1443 -5532
rect 1558 -5559 1575 -5532
rect 1690 -5559 1707 -5532
rect 1822 -5559 1839 -5532
rect 1954 -5559 1971 -5532
rect 1030 -5630 1047 -5603
rect 1030 -5630 1047 -5603
rect 1162 -5630 1179 -5603
rect 1294 -5630 1311 -5603
rect 1426 -5630 1443 -5603
rect 1558 -5630 1575 -5603
rect 1690 -5630 1707 -5603
rect 1822 -5630 1839 -5603
rect 1954 -5630 1971 -5603
rect 1030 -5701 1047 -5674
rect 1030 -5701 1047 -5674
rect 1162 -5701 1179 -5674
rect 1294 -5701 1311 -5674
rect 1426 -5701 1443 -5674
rect 1558 -5701 1575 -5674
rect 1690 -5701 1707 -5674
rect 1822 -5701 1839 -5674
rect 1954 -5701 1971 -5674
rect 1030 -5772 1047 -5745
rect 1030 -5772 1047 -5745
rect 1162 -5772 1179 -5745
rect 1294 -5772 1311 -5745
rect 1426 -5772 1443 -5745
rect 1558 -5772 1575 -5745
rect 1690 -5772 1707 -5745
rect 1822 -5772 1839 -5745
rect 1954 -5772 1971 -5745
rect 1030 -5843 1047 -5816
rect 1030 -5843 1047 -5816
rect 1162 -5843 1179 -5816
rect 1294 -5843 1311 -5816
rect 1426 -5843 1443 -5816
rect 1558 -5843 1575 -5816
rect 1690 -5843 1707 -5816
rect 1822 -5843 1839 -5816
rect 1954 -5843 1971 -5816
rect 1030 -5914 1047 -5887
rect 1030 -5914 1047 -5887
rect 1162 -5914 1179 -5887
rect 1294 -5914 1311 -5887
rect 1426 -5914 1443 -5887
rect 1558 -5914 1575 -5887
rect 1690 -5914 1707 -5887
rect 1822 -5914 1839 -5887
rect 1954 -5914 1971 -5887
rect 1030 -5985 1047 -5958
rect 1030 -5985 1047 -5958
rect 1162 -5985 1179 -5958
rect 1294 -5985 1311 -5958
rect 1426 -5985 1443 -5958
rect 1558 -5985 1575 -5958
rect 1690 -5985 1707 -5958
rect 1822 -5985 1839 -5958
rect 1954 -5985 1971 -5958
rect 1030 -6056 1047 -6029
rect 1030 -6056 1047 -6029
rect 1162 -6056 1179 -6029
rect 1294 -6056 1311 -6029
rect 1426 -6056 1443 -6029
rect 1558 -6056 1575 -6029
rect 1690 -6056 1707 -6029
rect 1822 -6056 1839 -6029
rect 1954 -6056 1971 -6029
rect 1030 -6127 1047 -6100
rect 1030 -6127 1047 -6100
rect 1162 -6127 1179 -6100
rect 1294 -6127 1311 -6100
rect 1426 -6127 1443 -6100
rect 1558 -6127 1575 -6100
rect 1690 -6127 1707 -6100
rect 1822 -6127 1839 -6100
rect 1954 -6127 1971 -6100
rect 1030 -6198 1047 -6171
rect 1030 -6198 1047 -6171
rect 1162 -6198 1179 -6171
rect 1294 -6198 1311 -6171
rect 1426 -6198 1443 -6171
rect 1558 -6198 1575 -6171
rect 1690 -6198 1707 -6171
rect 1822 -6198 1839 -6171
rect 1954 -6198 1971 -6171
rect 1030 -6269 1047 -6242
rect 1030 -6269 1047 -6242
rect 1162 -6269 1179 -6242
rect 1294 -6269 1311 -6242
rect 1426 -6269 1443 -6242
rect 1558 -6269 1575 -6242
rect 1690 -6269 1707 -6242
rect 1822 -6269 1839 -6242
rect 1954 -6269 1971 -6242
rect 1030 -6340 1047 -6313
rect 1030 -6340 1047 -6313
rect 1162 -6340 1179 -6313
rect 1294 -6340 1311 -6313
rect 1426 -6340 1443 -6313
rect 1558 -6340 1575 -6313
rect 1690 -6340 1707 -6313
rect 1822 -6340 1839 -6313
rect 1954 -6340 1971 -6313
rect 1030 -6411 1047 -6384
rect 1030 -6411 1047 -6384
rect 1162 -6411 1179 -6384
rect 1294 -6411 1311 -6384
rect 1426 -6411 1443 -6384
rect 1558 -6411 1575 -6384
rect 1690 -6411 1707 -6384
rect 1822 -6411 1839 -6384
rect 1954 -6411 1971 -6384
rect 1030 -6482 1047 -6455
rect 1030 -6482 1047 -6455
rect 1162 -6482 1179 -6455
rect 1294 -6482 1311 -6455
rect 1426 -6482 1443 -6455
rect 1558 -6482 1575 -6455
rect 1690 -6482 1707 -6455
rect 1822 -6482 1839 -6455
rect 1954 -6482 1971 -6455
rect 1030 -6553 1047 -6526
rect 1030 -6553 1047 -6526
rect 1162 -6553 1179 -6526
rect 1294 -6553 1311 -6526
rect 1426 -6553 1443 -6526
rect 1558 -6553 1575 -6526
rect 1690 -6553 1707 -6526
rect 1822 -6553 1839 -6526
rect 1954 -6553 1971 -6526
rect 1030 -6624 1047 -6597
rect 1030 -6624 1047 -6597
rect 1162 -6624 1179 -6597
rect 1294 -6624 1311 -6597
rect 1426 -6624 1443 -6597
rect 1558 -6624 1575 -6597
rect 1690 -6624 1707 -6597
rect 1822 -6624 1839 -6597
rect 1954 -6624 1971 -6597
rect 1030 -6695 1047 -6668
rect 1030 -6695 1047 -6668
rect 1162 -6695 1179 -6668
rect 1294 -6695 1311 -6668
rect 1426 -6695 1443 -6668
rect 1558 -6695 1575 -6668
rect 1690 -6695 1707 -6668
rect 1822 -6695 1839 -6668
rect 1954 -6695 1971 -6668
rect 1030 -6766 1047 -6739
rect 1030 -6766 1047 -6739
rect 1162 -6766 1179 -6739
rect 1294 -6766 1311 -6739
rect 1426 -6766 1443 -6739
rect 1558 -6766 1575 -6739
rect 1690 -6766 1707 -6739
rect 1822 -6766 1839 -6739
rect 1954 -6766 1971 -6739
rect 1030 -6837 1047 -6810
rect 1030 -6837 1047 -6810
rect 1162 -6837 1179 -6810
rect 1294 -6837 1311 -6810
rect 1426 -6837 1443 -6810
rect 1558 -6837 1575 -6810
rect 1690 -6837 1707 -6810
rect 1822 -6837 1839 -6810
rect 1954 -6837 1971 -6810
rect 1030 -6908 1047 -6881
rect 1030 -6908 1047 -6881
rect 1162 -6908 1179 -6881
rect 1294 -6908 1311 -6881
rect 1426 -6908 1443 -6881
rect 1558 -6908 1575 -6881
rect 1690 -6908 1707 -6881
rect 1822 -6908 1839 -6881
rect 1954 -6908 1971 -6881
rect 1030 -6979 1047 -6952
rect 1030 -6979 1047 -6952
rect 1162 -6979 1179 -6952
rect 1294 -6979 1311 -6952
rect 1426 -6979 1443 -6952
rect 1558 -6979 1575 -6952
rect 1690 -6979 1707 -6952
rect 1822 -6979 1839 -6952
rect 1954 -6979 1971 -6952
rect 1030 -7050 1047 -7023
rect 1030 -7050 1047 -7023
rect 1162 -7050 1179 -7023
rect 1294 -7050 1311 -7023
rect 1426 -7050 1443 -7023
rect 1558 -7050 1575 -7023
rect 1690 -7050 1707 -7023
rect 1822 -7050 1839 -7023
rect 1954 -7050 1971 -7023
rect 1030 -7121 1047 -7094
rect 1030 -7121 1047 -7094
rect 1162 -7121 1179 -7094
rect 1294 -7121 1311 -7094
rect 1426 -7121 1443 -7094
rect 1558 -7121 1575 -7094
rect 1690 -7121 1707 -7094
rect 1822 -7121 1839 -7094
rect 1954 -7121 1971 -7094
rect 1030 -7192 1047 -7165
rect 1030 -7192 1047 -7165
rect 1162 -7192 1179 -7165
rect 1294 -7192 1311 -7165
rect 1426 -7192 1443 -7165
rect 1558 -7192 1575 -7165
rect 1690 -7192 1707 -7165
rect 1822 -7192 1839 -7165
rect 1954 -7192 1971 -7165
rect 1030 -7263 1047 -7236
rect 1030 -7263 1047 -7236
rect 1162 -7263 1179 -7236
rect 1294 -7263 1311 -7236
rect 1426 -7263 1443 -7236
rect 1558 -7263 1575 -7236
rect 1690 -7263 1707 -7236
rect 1822 -7263 1839 -7236
rect 1954 -7263 1971 -7236
rect 1030 -7334 1047 -7307
rect 1030 -7334 1047 -7307
rect 1162 -7334 1179 -7307
rect 1294 -7334 1311 -7307
rect 1426 -7334 1443 -7307
rect 1558 -7334 1575 -7307
rect 1690 -7334 1707 -7307
rect 1822 -7334 1839 -7307
rect 1954 -7334 1971 -7307
rect 1030 -7405 1047 -7378
rect 1030 -7405 1047 -7378
rect 1162 -7405 1179 -7378
rect 1294 -7405 1311 -7378
rect 1426 -7405 1443 -7378
rect 1558 -7405 1575 -7378
rect 1690 -7405 1707 -7378
rect 1822 -7405 1839 -7378
rect 1954 -7405 1971 -7378
rect 1030 -7476 1047 -7449
rect 1030 -7476 1047 -7449
rect 1162 -7476 1179 -7449
rect 1294 -7476 1311 -7449
rect 1426 -7476 1443 -7449
rect 1558 -7476 1575 -7449
rect 1690 -7476 1707 -7449
rect 1822 -7476 1839 -7449
rect 1954 -7476 1971 -7449
rect 1030 -7547 1047 -7520
rect 1030 -7547 1047 -7520
rect 1162 -7547 1179 -7520
rect 1294 -7547 1311 -7520
rect 1426 -7547 1443 -7520
rect 1558 -7547 1575 -7520
rect 1690 -7547 1707 -7520
rect 1822 -7547 1839 -7520
rect 1954 -7547 1971 -7520
rect 1030 -7618 1047 -7591
rect 1030 -7618 1047 -7591
rect 1162 -7618 1179 -7591
rect 1294 -7618 1311 -7591
rect 1426 -7618 1443 -7591
rect 1558 -7618 1575 -7591
rect 1690 -7618 1707 -7591
rect 1822 -7618 1839 -7591
rect 1954 -7618 1971 -7591
rect 1030 -7689 1047 -7662
rect 1030 -7689 1047 -7662
rect 1162 -7689 1179 -7662
rect 1294 -7689 1311 -7662
rect 1426 -7689 1443 -7662
rect 1558 -7689 1575 -7662
rect 1690 -7689 1707 -7662
rect 1822 -7689 1839 -7662
rect 1954 -7689 1971 -7662
rect 1030 -7760 1047 -7733
rect 1030 -7760 1047 -7733
rect 1162 -7760 1179 -7733
rect 1294 -7760 1311 -7733
rect 1426 -7760 1443 -7733
rect 1558 -7760 1575 -7733
rect 1690 -7760 1707 -7733
rect 1822 -7760 1839 -7733
rect 1954 -7760 1971 -7733
rect 1030 -7831 1047 -7804
rect 1030 -7831 1047 -7804
rect 1162 -7831 1179 -7804
rect 1294 -7831 1311 -7804
rect 1426 -7831 1443 -7804
rect 1558 -7831 1575 -7804
rect 1690 -7831 1707 -7804
rect 1822 -7831 1839 -7804
rect 1954 -7831 1971 -7804
rect 1030 -7902 1047 -7875
rect 1030 -7902 1047 -7875
rect 1162 -7902 1179 -7875
rect 1294 -7902 1311 -7875
rect 1426 -7902 1443 -7875
rect 1558 -7902 1575 -7875
rect 1690 -7902 1707 -7875
rect 1822 -7902 1839 -7875
rect 1954 -7902 1971 -7875
rect 1030 -7973 1047 -7946
rect 1030 -7973 1047 -7946
rect 1162 -7973 1179 -7946
rect 1294 -7973 1311 -7946
rect 1426 -7973 1443 -7946
rect 1558 -7973 1575 -7946
rect 1690 -7973 1707 -7946
rect 1822 -7973 1839 -7946
rect 1954 -7973 1971 -7946
rect 1030 -8044 1047 -8017
rect 1030 -8044 1047 -8017
rect 1162 -8044 1179 -8017
rect 1294 -8044 1311 -8017
rect 1426 -8044 1443 -8017
rect 1558 -8044 1575 -8017
rect 1690 -8044 1707 -8017
rect 1822 -8044 1839 -8017
rect 1954 -8044 1971 -8017
rect 1030 -8115 1047 -8088
rect 1030 -8115 1047 -8088
rect 1162 -8115 1179 -8088
rect 1294 -8115 1311 -8088
rect 1426 -8115 1443 -8088
rect 1558 -8115 1575 -8088
rect 1690 -8115 1707 -8088
rect 1822 -8115 1839 -8088
rect 1954 -8115 1971 -8088
rect 1030 -8186 1047 -8159
rect 1030 -8186 1047 -8159
rect 1162 -8186 1179 -8159
rect 1294 -8186 1311 -8159
rect 1426 -8186 1443 -8159
rect 1558 -8186 1575 -8159
rect 1690 -8186 1707 -8159
rect 1822 -8186 1839 -8159
rect 1954 -8186 1971 -8159
rect 1030 -8257 1047 -8230
rect 1030 -8257 1047 -8230
rect 1162 -8257 1179 -8230
rect 1294 -8257 1311 -8230
rect 1426 -8257 1443 -8230
rect 1558 -8257 1575 -8230
rect 1690 -8257 1707 -8230
rect 1822 -8257 1839 -8230
rect 1954 -8257 1971 -8230
rect 1030 -8328 1047 -8301
rect 1030 -8328 1047 -8301
rect 1162 -8328 1179 -8301
rect 1294 -8328 1311 -8301
rect 1426 -8328 1443 -8301
rect 1558 -8328 1575 -8301
rect 1690 -8328 1707 -8301
rect 1822 -8328 1839 -8301
rect 1954 -8328 1971 -8301
rect 1030 -8399 1047 -8372
rect 1030 -8399 1047 -8372
rect 1162 -8399 1179 -8372
rect 1294 -8399 1311 -8372
rect 1426 -8399 1443 -8372
rect 1558 -8399 1575 -8372
rect 1690 -8399 1707 -8372
rect 1822 -8399 1839 -8372
rect 1954 -8399 1971 -8372
rect 1030 -8470 1047 -8443
rect 1030 -8470 1047 -8443
rect 1162 -8470 1179 -8443
rect 1294 -8470 1311 -8443
rect 1426 -8470 1443 -8443
rect 1558 -8470 1575 -8443
rect 1690 -8470 1707 -8443
rect 1822 -8470 1839 -8443
rect 1954 -8470 1971 -8443
rect 1030 -8541 1047 -8514
rect 1030 -8541 1047 -8514
rect 1162 -8541 1179 -8514
rect 1294 -8541 1311 -8514
rect 1426 -8541 1443 -8514
rect 1558 -8541 1575 -8514
rect 1690 -8541 1707 -8514
rect 1822 -8541 1839 -8514
rect 1954 -8541 1971 -8514
rect 1030 -8612 1047 -8585
rect 1030 -8612 1047 -8585
rect 1162 -8612 1179 -8585
rect 1294 -8612 1311 -8585
rect 1426 -8612 1443 -8585
rect 1558 -8612 1575 -8585
rect 1690 -8612 1707 -8585
rect 1822 -8612 1839 -8585
rect 1954 -8612 1971 -8585
rect 1030 -8683 1047 -8656
rect 1030 -8683 1047 -8656
rect 1162 -8683 1179 -8656
rect 1294 -8683 1311 -8656
rect 1426 -8683 1443 -8656
rect 1558 -8683 1575 -8656
rect 1690 -8683 1707 -8656
rect 1822 -8683 1839 -8656
rect 1954 -8683 1971 -8656
rect 1030 -8754 1047 -8727
rect 1030 -8754 1047 -8727
rect 1162 -8754 1179 -8727
rect 1294 -8754 1311 -8727
rect 1426 -8754 1443 -8727
rect 1558 -8754 1575 -8727
rect 1690 -8754 1707 -8727
rect 1822 -8754 1839 -8727
rect 1954 -8754 1971 -8727
rect 1030 -8825 1047 -8798
rect 1030 -8825 1047 -8798
rect 1162 -8825 1179 -8798
rect 1294 -8825 1311 -8798
rect 1426 -8825 1443 -8798
rect 1558 -8825 1575 -8798
rect 1690 -8825 1707 -8798
rect 1822 -8825 1839 -8798
rect 1954 -8825 1971 -8798
rect 1030 -8896 1047 -8869
rect 1030 -8896 1047 -8869
rect 1162 -8896 1179 -8869
rect 1294 -8896 1311 -8869
rect 1426 -8896 1443 -8869
rect 1558 -8896 1575 -8869
rect 1690 -8896 1707 -8869
rect 1822 -8896 1839 -8869
rect 1954 -8896 1971 -8869
rect 1030 -8967 1047 -8940
rect 1030 -8967 1047 -8940
rect 1162 -8967 1179 -8940
rect 1294 -8967 1311 -8940
rect 1426 -8967 1443 -8940
rect 1558 -8967 1575 -8940
rect 1690 -8967 1707 -8940
rect 1822 -8967 1839 -8940
rect 1954 -8967 1971 -8940
rect 1030 -9038 1047 -9011
rect 1030 -9038 1047 -9011
rect 1162 -9038 1179 -9011
rect 1294 -9038 1311 -9011
rect 1426 -9038 1443 -9011
rect 1558 -9038 1575 -9011
rect 1690 -9038 1707 -9011
rect 1822 -9038 1839 -9011
rect 1954 -9038 1971 -9011
rect 1030 -9109 1047 -9082
rect 1030 -9109 1047 -9082
rect 1162 -9109 1179 -9082
rect 1294 -9109 1311 -9082
rect 1426 -9109 1443 -9082
rect 1558 -9109 1575 -9082
rect 1690 -9109 1707 -9082
rect 1822 -9109 1839 -9082
rect 1954 -9109 1971 -9082
rect 8 90 25 117
rect 64 150 81 167
rect 140 90 157 117
rect 196 150 213 167
rect 272 90 289 117
rect 328 150 345 167
rect 404 90 421 117
rect 460 150 477 167
rect 536 90 553 117
rect 592 150 609 167
rect 668 90 685 117
rect 724 150 741 167
rect 800 90 817 117
rect 856 150 873 167
rect 1129 90 1146 117
rect 1073 150 1090 167
rect 1261 90 1278 117
rect 1205 150 1222 167
rect 1393 90 1410 117
rect 1337 150 1354 167
rect 1525 90 1542 117
rect 1469 150 1486 167
rect 1657 90 1674 117
rect 1601 150 1618 167
rect 1789 90 1806 117
rect 1733 150 1750 167
rect 1921 90 1938 117
rect 1865 150 1882 167
<< metal1 >>
rect 0 -33 33 0
rect 66 -33 99 0
rect 132 -33 165 0
rect 198 -33 231 0
rect 264 -33 297 0
rect 330 -33 363 0
rect 396 -33 429 0
rect 462 -33 495 0
rect 528 -33 561 0
rect 594 -33 627 0
rect 660 -33 693 0
rect 726 -33 759 0
rect 792 -33 825 0
rect 858 -33 891 0
rect 1055 -33 1088 0
rect 1121 -33 1154 0
rect 1187 -33 1220 0
rect 1253 -33 1286 0
rect 1319 -33 1352 0
rect 1385 -33 1418 0
rect 1451 -33 1484 0
rect 1517 -33 1550 0
rect 1583 -33 1616 0
rect 1649 -33 1682 0
rect 1715 -33 1748 0
rect 1781 -33 1814 0
rect 1847 -33 1880 0
rect 1913 -33 1946 0
rect 1022 -100 1979 -57
rect 1022 -171 1979 -128
rect 1022 -242 1979 -199
rect 1022 -313 1979 -270
rect 1022 -384 1979 -341
rect 1022 -455 1979 -412
rect 1022 -526 1979 -483
rect 1022 -597 1979 -554
rect 1022 -668 1979 -625
rect 1022 -739 1979 -696
rect 1022 -810 1979 -767
rect 1022 -881 1979 -838
rect 1022 -952 1979 -909
rect 1022 -1023 1979 -980
rect 1022 -1094 1979 -1051
rect 1022 -1165 1979 -1122
rect 1022 -1236 1979 -1193
rect 1022 -1307 1979 -1264
rect 1022 -1378 1979 -1335
rect 1022 -1449 1979 -1406
rect 1022 -1520 1979 -1477
rect 1022 -1591 1979 -1548
rect 1022 -1662 1979 -1619
rect 1022 -1733 1979 -1690
rect 1022 -1804 1979 -1761
rect 1022 -1875 1979 -1832
rect 1022 -1946 1979 -1903
rect 1022 -2017 1979 -1974
rect 1022 -2088 1979 -2045
rect 1022 -2159 1979 -2116
rect 1022 -2230 1979 -2187
rect 1022 -2301 1979 -2258
rect 1022 -2372 1979 -2329
rect 1022 -2443 1979 -2400
rect 1022 -2514 1979 -2471
rect 1022 -2585 1979 -2542
rect 1022 -2656 1979 -2613
rect 1022 -2727 1979 -2684
rect 1022 -2798 1979 -2755
rect 1022 -2869 1979 -2826
rect 1022 -2940 1979 -2897
rect 1022 -3011 1979 -2968
rect 1022 -3082 1979 -3039
rect 1022 -3153 1979 -3110
rect 1022 -3224 1979 -3181
rect 1022 -3295 1979 -3252
rect 1022 -3366 1979 -3323
rect 1022 -3437 1979 -3394
rect 1022 -3508 1979 -3465
rect 1022 -3579 1979 -3536
rect 1022 -3650 1979 -3607
rect 1022 -3721 1979 -3678
rect 1022 -3792 1979 -3749
rect 1022 -3863 1979 -3820
rect 1022 -3934 1979 -3891
rect 1022 -4005 1979 -3962
rect 1022 -4076 1979 -4033
rect 1022 -4147 1979 -4104
rect 1022 -4218 1979 -4175
rect 1022 -4289 1979 -4246
rect 1022 -4360 1979 -4317
rect 1022 -4431 1979 -4388
rect 1022 -4502 1979 -4459
rect 1022 -4573 1979 -4530
rect 1022 -4644 1979 -4601
rect 1022 -4715 1979 -4672
rect 1022 -4786 1979 -4743
rect 1022 -4857 1979 -4814
rect 1022 -4928 1979 -4885
rect 1022 -4999 1979 -4956
rect 1022 -5070 1979 -5027
rect 1022 -5141 1979 -5098
rect 1022 -5212 1979 -5169
rect 1022 -5283 1979 -5240
rect 1022 -5354 1979 -5311
rect 1022 -5425 1979 -5382
rect 1022 -5496 1979 -5453
rect 1022 -5567 1979 -5524
rect 1022 -5638 1979 -5595
rect 1022 -5709 1979 -5666
rect 1022 -5780 1979 -5737
rect 1022 -5851 1979 -5808
rect 1022 -5922 1979 -5879
rect 1022 -5993 1979 -5950
rect 1022 -6064 1979 -6021
rect 1022 -6135 1979 -6092
rect 1022 -6206 1979 -6163
rect 1022 -6277 1979 -6234
rect 1022 -6348 1979 -6305
rect 1022 -6419 1979 -6376
rect 1022 -6490 1979 -6447
rect 1022 -6561 1979 -6518
rect 1022 -6632 1979 -6589
rect 1022 -6703 1979 -6660
rect 1022 -6774 1979 -6731
rect 1022 -6845 1979 -6802
rect 1022 -6916 1979 -6873
rect 1022 -6987 1979 -6944
rect 1022 -7058 1979 -7015
rect 1022 -7129 1979 -7086
rect 1022 -7200 1979 -7157
rect 1022 -7271 1979 -7228
rect 1022 -7342 1979 -7299
rect 1022 -7413 1979 -7370
rect 1022 -7484 1979 -7441
rect 1022 -7555 1979 -7512
rect 1022 -7626 1979 -7583
rect 1022 -7697 1979 -7654
rect 1022 -7768 1979 -7725
rect 1022 -7839 1979 -7796
rect 1022 -7910 1979 -7867
rect 1022 -7981 1979 -7938
rect 1022 -8052 1979 -8009
rect 1022 -8123 1979 -8080
rect 1022 -8194 1979 -8151
rect 1022 -8265 1979 -8222
rect 1022 -8336 1979 -8293
rect 1022 -8407 1979 -8364
rect 1022 -8478 1979 -8435
rect 1022 -8549 1979 -8506
rect 1022 -8620 1979 -8577
rect 1022 -8691 1979 -8648
rect 1022 -8762 1979 -8719
rect 1022 -8833 1979 -8790
rect 1022 -8904 1979 -8861
rect 1022 -8975 1979 -8932
rect 1022 -9046 1979 -9003
rect 1022 -9117 1979 -9074
rect 0 0 33 125
rect 56 142 89 175
rect 66 0 99 175
rect 132 0 165 125
rect 188 142 221 175
rect 198 0 231 175
rect 264 0 297 125
rect 320 142 353 175
rect 330 0 363 175
rect 396 0 429 125
rect 452 142 485 175
rect 462 0 495 175
rect 528 0 561 125
rect 584 142 617 175
rect 594 0 627 175
rect 660 0 693 125
rect 716 142 749 175
rect 726 0 759 175
rect 792 0 825 125
rect 848 142 881 175
rect 858 0 891 175
rect 858 175 891 175
rect 1055 175 1088 175
rect 891 142 1055 175
rect 726 175 759 222
rect 1187 175 1220 222
rect 759 189 1187 222
rect 594 175 627 269
rect 1319 175 1352 269
rect 627 236 1319 269
rect 462 175 495 316
rect 1451 175 1484 316
rect 495 283 1451 316
rect 330 175 363 363
rect 1583 175 1616 363
rect 363 330 1583 363
rect 198 175 231 410
rect 1715 175 1748 410
rect 231 377 1715 410
rect 66 175 99 457
rect 1847 175 1880 457
rect 99 424 1847 457
rect 1121 0 1154 125
rect 1065 142 1098 175
rect 1055 0 1088 175
rect 1253 0 1286 125
rect 1197 142 1230 175
rect 1187 0 1220 175
rect 1385 0 1418 125
rect 1329 142 1362 175
rect 1319 0 1352 175
rect 1517 0 1550 125
rect 1461 142 1494 175
rect 1451 0 1484 175
rect 1649 0 1682 125
rect 1593 142 1626 175
rect 1583 0 1616 175
rect 1781 0 1814 125
rect 1725 142 1758 175
rect 1715 0 1748 175
rect 1913 0 1946 125
rect 1857 142 1890 175
rect 1847 0 1880 175
<< via1 >>
rect 894 145 921 172
rect 762 192 789 219
rect 630 239 657 266
rect 498 286 525 313
rect 366 333 393 360
rect 234 380 261 407
rect 102 427 129 454
<< metal2 >>
rect 891 142 924 175
rect 759 189 792 222
rect 627 236 660 269
rect 495 283 528 316
rect 363 330 396 363
rect 231 377 264 410
rect 99 424 132 457
<< pdiff >>
rect -33 -100 0 -57
rect 33 -100 66 -57
rect 66 -100 99 -57
rect 99 -100 132 -57
rect 165 -100 198 -57
rect 198 -100 231 -57
rect 231 -100 264 -57
rect 297 -100 330 -57
rect 330 -100 363 -57
rect 363 -100 396 -57
rect 429 -100 462 -57
rect 462 -100 495 -57
rect 495 -100 528 -57
rect 561 -100 594 -57
rect 594 -100 627 -57
rect 627 -100 660 -57
rect 693 -100 726 -57
rect 726 -100 759 -57
rect 759 -100 792 -57
rect 825 -100 858 -57
rect 858 -100 891 -57
rect 891 -100 924 -57
rect -33 -171 0 -128
rect 33 -171 66 -128
rect 66 -171 99 -128
rect 99 -171 132 -128
rect 165 -171 198 -128
rect 198 -171 231 -128
rect 231 -171 264 -128
rect 297 -171 330 -128
rect 330 -171 363 -128
rect 363 -171 396 -128
rect 429 -171 462 -128
rect 462 -171 495 -128
rect 495 -171 528 -128
rect 561 -171 594 -128
rect 594 -171 627 -128
rect 627 -171 660 -128
rect 693 -171 726 -128
rect 726 -171 759 -128
rect 759 -171 792 -128
rect 825 -171 858 -128
rect 792 -171 825 -128
rect 891 -171 924 -128
rect -33 -242 0 -199
rect 33 -242 66 -199
rect 66 -242 99 -199
rect 99 -242 132 -199
rect 165 -242 198 -199
rect 198 -242 231 -199
rect 231 -242 264 -199
rect 297 -242 330 -199
rect 330 -242 363 -199
rect 363 -242 396 -199
rect 429 -242 462 -199
rect 462 -242 495 -199
rect 495 -242 528 -199
rect 561 -242 594 -199
rect 594 -242 627 -199
rect 627 -242 660 -199
rect 693 -242 726 -199
rect 660 -242 693 -199
rect 759 -242 792 -199
rect 825 -242 858 -199
rect 858 -242 891 -199
rect 891 -242 924 -199
rect -33 -313 0 -270
rect 33 -313 66 -270
rect 66 -313 99 -270
rect 99 -313 132 -270
rect 165 -313 198 -270
rect 198 -313 231 -270
rect 231 -313 264 -270
rect 297 -313 330 -270
rect 330 -313 363 -270
rect 363 -313 396 -270
rect 429 -313 462 -270
rect 462 -313 495 -270
rect 495 -313 528 -270
rect 561 -313 594 -270
rect 594 -313 627 -270
rect 627 -313 660 -270
rect 693 -313 726 -270
rect 660 -313 693 -270
rect 759 -313 792 -270
rect 825 -313 858 -270
rect 792 -313 825 -270
rect 891 -313 924 -270
rect -33 -384 0 -341
rect 33 -384 66 -341
rect 66 -384 99 -341
rect 99 -384 132 -341
rect 165 -384 198 -341
rect 198 -384 231 -341
rect 231 -384 264 -341
rect 297 -384 330 -341
rect 330 -384 363 -341
rect 363 -384 396 -341
rect 429 -384 462 -341
rect 462 -384 495 -341
rect 495 -384 528 -341
rect 561 -384 594 -341
rect 528 -384 561 -341
rect 627 -384 660 -341
rect 693 -384 726 -341
rect 726 -384 759 -341
rect 759 -384 792 -341
rect 825 -384 858 -341
rect 858 -384 891 -341
rect 891 -384 924 -341
rect -33 -455 0 -412
rect 33 -455 66 -412
rect 66 -455 99 -412
rect 99 -455 132 -412
rect 165 -455 198 -412
rect 198 -455 231 -412
rect 231 -455 264 -412
rect 297 -455 330 -412
rect 330 -455 363 -412
rect 363 -455 396 -412
rect 429 -455 462 -412
rect 462 -455 495 -412
rect 495 -455 528 -412
rect 561 -455 594 -412
rect 528 -455 561 -412
rect 627 -455 660 -412
rect 693 -455 726 -412
rect 726 -455 759 -412
rect 759 -455 792 -412
rect 825 -455 858 -412
rect 792 -455 825 -412
rect 891 -455 924 -412
rect -33 -526 0 -483
rect 33 -526 66 -483
rect 66 -526 99 -483
rect 99 -526 132 -483
rect 165 -526 198 -483
rect 198 -526 231 -483
rect 231 -526 264 -483
rect 297 -526 330 -483
rect 330 -526 363 -483
rect 363 -526 396 -483
rect 429 -526 462 -483
rect 462 -526 495 -483
rect 495 -526 528 -483
rect 561 -526 594 -483
rect 528 -526 561 -483
rect 627 -526 660 -483
rect 693 -526 726 -483
rect 660 -526 693 -483
rect 759 -526 792 -483
rect 825 -526 858 -483
rect 858 -526 891 -483
rect 891 -526 924 -483
rect -33 -597 0 -554
rect 33 -597 66 -554
rect 66 -597 99 -554
rect 99 -597 132 -554
rect 165 -597 198 -554
rect 198 -597 231 -554
rect 231 -597 264 -554
rect 297 -597 330 -554
rect 330 -597 363 -554
rect 363 -597 396 -554
rect 429 -597 462 -554
rect 462 -597 495 -554
rect 495 -597 528 -554
rect 561 -597 594 -554
rect 528 -597 561 -554
rect 627 -597 660 -554
rect 693 -597 726 -554
rect 660 -597 693 -554
rect 759 -597 792 -554
rect 825 -597 858 -554
rect 792 -597 825 -554
rect 891 -597 924 -554
rect -33 -668 0 -625
rect 33 -668 66 -625
rect 66 -668 99 -625
rect 99 -668 132 -625
rect 165 -668 198 -625
rect 198 -668 231 -625
rect 231 -668 264 -625
rect 297 -668 330 -625
rect 330 -668 363 -625
rect 363 -668 396 -625
rect 429 -668 462 -625
rect 396 -668 429 -625
rect 495 -668 528 -625
rect 561 -668 594 -625
rect 594 -668 627 -625
rect 627 -668 660 -625
rect 693 -668 726 -625
rect 726 -668 759 -625
rect 759 -668 792 -625
rect 825 -668 858 -625
rect 858 -668 891 -625
rect 891 -668 924 -625
rect -33 -739 0 -696
rect 33 -739 66 -696
rect 66 -739 99 -696
rect 99 -739 132 -696
rect 165 -739 198 -696
rect 198 -739 231 -696
rect 231 -739 264 -696
rect 297 -739 330 -696
rect 330 -739 363 -696
rect 363 -739 396 -696
rect 429 -739 462 -696
rect 396 -739 429 -696
rect 495 -739 528 -696
rect 561 -739 594 -696
rect 594 -739 627 -696
rect 627 -739 660 -696
rect 693 -739 726 -696
rect 726 -739 759 -696
rect 759 -739 792 -696
rect 825 -739 858 -696
rect 792 -739 825 -696
rect 891 -739 924 -696
rect -33 -810 0 -767
rect 33 -810 66 -767
rect 66 -810 99 -767
rect 99 -810 132 -767
rect 165 -810 198 -767
rect 198 -810 231 -767
rect 231 -810 264 -767
rect 297 -810 330 -767
rect 330 -810 363 -767
rect 363 -810 396 -767
rect 429 -810 462 -767
rect 396 -810 429 -767
rect 495 -810 528 -767
rect 561 -810 594 -767
rect 594 -810 627 -767
rect 627 -810 660 -767
rect 693 -810 726 -767
rect 660 -810 693 -767
rect 759 -810 792 -767
rect 825 -810 858 -767
rect 858 -810 891 -767
rect 891 -810 924 -767
rect -33 -881 0 -838
rect 33 -881 66 -838
rect 66 -881 99 -838
rect 99 -881 132 -838
rect 165 -881 198 -838
rect 198 -881 231 -838
rect 231 -881 264 -838
rect 297 -881 330 -838
rect 330 -881 363 -838
rect 363 -881 396 -838
rect 429 -881 462 -838
rect 396 -881 429 -838
rect 495 -881 528 -838
rect 561 -881 594 -838
rect 594 -881 627 -838
rect 627 -881 660 -838
rect 693 -881 726 -838
rect 660 -881 693 -838
rect 759 -881 792 -838
rect 825 -881 858 -838
rect 792 -881 825 -838
rect 891 -881 924 -838
rect -33 -952 0 -909
rect 33 -952 66 -909
rect 66 -952 99 -909
rect 99 -952 132 -909
rect 165 -952 198 -909
rect 198 -952 231 -909
rect 231 -952 264 -909
rect 297 -952 330 -909
rect 330 -952 363 -909
rect 363 -952 396 -909
rect 429 -952 462 -909
rect 396 -952 429 -909
rect 495 -952 528 -909
rect 561 -952 594 -909
rect 528 -952 561 -909
rect 627 -952 660 -909
rect 693 -952 726 -909
rect 726 -952 759 -909
rect 759 -952 792 -909
rect 825 -952 858 -909
rect 858 -952 891 -909
rect 891 -952 924 -909
rect -33 -1023 0 -980
rect 33 -1023 66 -980
rect 66 -1023 99 -980
rect 99 -1023 132 -980
rect 165 -1023 198 -980
rect 198 -1023 231 -980
rect 231 -1023 264 -980
rect 297 -1023 330 -980
rect 330 -1023 363 -980
rect 363 -1023 396 -980
rect 429 -1023 462 -980
rect 396 -1023 429 -980
rect 495 -1023 528 -980
rect 561 -1023 594 -980
rect 528 -1023 561 -980
rect 627 -1023 660 -980
rect 693 -1023 726 -980
rect 726 -1023 759 -980
rect 759 -1023 792 -980
rect 825 -1023 858 -980
rect 792 -1023 825 -980
rect 891 -1023 924 -980
rect -33 -1094 0 -1051
rect 33 -1094 66 -1051
rect 66 -1094 99 -1051
rect 99 -1094 132 -1051
rect 165 -1094 198 -1051
rect 198 -1094 231 -1051
rect 231 -1094 264 -1051
rect 297 -1094 330 -1051
rect 330 -1094 363 -1051
rect 363 -1094 396 -1051
rect 429 -1094 462 -1051
rect 396 -1094 429 -1051
rect 495 -1094 528 -1051
rect 561 -1094 594 -1051
rect 528 -1094 561 -1051
rect 627 -1094 660 -1051
rect 693 -1094 726 -1051
rect 660 -1094 693 -1051
rect 759 -1094 792 -1051
rect 825 -1094 858 -1051
rect 858 -1094 891 -1051
rect 891 -1094 924 -1051
rect -33 -1165 0 -1122
rect 33 -1165 66 -1122
rect 66 -1165 99 -1122
rect 99 -1165 132 -1122
rect 165 -1165 198 -1122
rect 198 -1165 231 -1122
rect 231 -1165 264 -1122
rect 297 -1165 330 -1122
rect 330 -1165 363 -1122
rect 363 -1165 396 -1122
rect 429 -1165 462 -1122
rect 396 -1165 429 -1122
rect 495 -1165 528 -1122
rect 561 -1165 594 -1122
rect 528 -1165 561 -1122
rect 627 -1165 660 -1122
rect 693 -1165 726 -1122
rect 660 -1165 693 -1122
rect 759 -1165 792 -1122
rect 825 -1165 858 -1122
rect 792 -1165 825 -1122
rect 891 -1165 924 -1122
rect -33 -1236 0 -1193
rect 33 -1236 66 -1193
rect 66 -1236 99 -1193
rect 99 -1236 132 -1193
rect 165 -1236 198 -1193
rect 198 -1236 231 -1193
rect 231 -1236 264 -1193
rect 297 -1236 330 -1193
rect 264 -1236 297 -1193
rect 363 -1236 396 -1193
rect 429 -1236 462 -1193
rect 462 -1236 495 -1193
rect 495 -1236 528 -1193
rect 561 -1236 594 -1193
rect 594 -1236 627 -1193
rect 627 -1236 660 -1193
rect 693 -1236 726 -1193
rect 726 -1236 759 -1193
rect 759 -1236 792 -1193
rect 825 -1236 858 -1193
rect 858 -1236 891 -1193
rect 891 -1236 924 -1193
rect -33 -1307 0 -1264
rect 33 -1307 66 -1264
rect 66 -1307 99 -1264
rect 99 -1307 132 -1264
rect 165 -1307 198 -1264
rect 198 -1307 231 -1264
rect 231 -1307 264 -1264
rect 297 -1307 330 -1264
rect 264 -1307 297 -1264
rect 363 -1307 396 -1264
rect 429 -1307 462 -1264
rect 462 -1307 495 -1264
rect 495 -1307 528 -1264
rect 561 -1307 594 -1264
rect 594 -1307 627 -1264
rect 627 -1307 660 -1264
rect 693 -1307 726 -1264
rect 726 -1307 759 -1264
rect 759 -1307 792 -1264
rect 825 -1307 858 -1264
rect 792 -1307 825 -1264
rect 891 -1307 924 -1264
rect -33 -1378 0 -1335
rect 33 -1378 66 -1335
rect 66 -1378 99 -1335
rect 99 -1378 132 -1335
rect 165 -1378 198 -1335
rect 198 -1378 231 -1335
rect 231 -1378 264 -1335
rect 297 -1378 330 -1335
rect 264 -1378 297 -1335
rect 363 -1378 396 -1335
rect 429 -1378 462 -1335
rect 462 -1378 495 -1335
rect 495 -1378 528 -1335
rect 561 -1378 594 -1335
rect 594 -1378 627 -1335
rect 627 -1378 660 -1335
rect 693 -1378 726 -1335
rect 660 -1378 693 -1335
rect 759 -1378 792 -1335
rect 825 -1378 858 -1335
rect 858 -1378 891 -1335
rect 891 -1378 924 -1335
rect -33 -1449 0 -1406
rect 33 -1449 66 -1406
rect 66 -1449 99 -1406
rect 99 -1449 132 -1406
rect 165 -1449 198 -1406
rect 198 -1449 231 -1406
rect 231 -1449 264 -1406
rect 297 -1449 330 -1406
rect 264 -1449 297 -1406
rect 363 -1449 396 -1406
rect 429 -1449 462 -1406
rect 462 -1449 495 -1406
rect 495 -1449 528 -1406
rect 561 -1449 594 -1406
rect 594 -1449 627 -1406
rect 627 -1449 660 -1406
rect 693 -1449 726 -1406
rect 660 -1449 693 -1406
rect 759 -1449 792 -1406
rect 825 -1449 858 -1406
rect 792 -1449 825 -1406
rect 891 -1449 924 -1406
rect -33 -1520 0 -1477
rect 33 -1520 66 -1477
rect 66 -1520 99 -1477
rect 99 -1520 132 -1477
rect 165 -1520 198 -1477
rect 198 -1520 231 -1477
rect 231 -1520 264 -1477
rect 297 -1520 330 -1477
rect 264 -1520 297 -1477
rect 363 -1520 396 -1477
rect 429 -1520 462 -1477
rect 462 -1520 495 -1477
rect 495 -1520 528 -1477
rect 561 -1520 594 -1477
rect 528 -1520 561 -1477
rect 627 -1520 660 -1477
rect 693 -1520 726 -1477
rect 726 -1520 759 -1477
rect 759 -1520 792 -1477
rect 825 -1520 858 -1477
rect 858 -1520 891 -1477
rect 891 -1520 924 -1477
rect -33 -1591 0 -1548
rect 33 -1591 66 -1548
rect 66 -1591 99 -1548
rect 99 -1591 132 -1548
rect 165 -1591 198 -1548
rect 198 -1591 231 -1548
rect 231 -1591 264 -1548
rect 297 -1591 330 -1548
rect 264 -1591 297 -1548
rect 363 -1591 396 -1548
rect 429 -1591 462 -1548
rect 462 -1591 495 -1548
rect 495 -1591 528 -1548
rect 561 -1591 594 -1548
rect 528 -1591 561 -1548
rect 627 -1591 660 -1548
rect 693 -1591 726 -1548
rect 726 -1591 759 -1548
rect 759 -1591 792 -1548
rect 825 -1591 858 -1548
rect 792 -1591 825 -1548
rect 891 -1591 924 -1548
rect -33 -1662 0 -1619
rect 33 -1662 66 -1619
rect 66 -1662 99 -1619
rect 99 -1662 132 -1619
rect 165 -1662 198 -1619
rect 198 -1662 231 -1619
rect 231 -1662 264 -1619
rect 297 -1662 330 -1619
rect 264 -1662 297 -1619
rect 363 -1662 396 -1619
rect 429 -1662 462 -1619
rect 462 -1662 495 -1619
rect 495 -1662 528 -1619
rect 561 -1662 594 -1619
rect 528 -1662 561 -1619
rect 627 -1662 660 -1619
rect 693 -1662 726 -1619
rect 660 -1662 693 -1619
rect 759 -1662 792 -1619
rect 825 -1662 858 -1619
rect 858 -1662 891 -1619
rect 891 -1662 924 -1619
rect -33 -1733 0 -1690
rect 33 -1733 66 -1690
rect 66 -1733 99 -1690
rect 99 -1733 132 -1690
rect 165 -1733 198 -1690
rect 198 -1733 231 -1690
rect 231 -1733 264 -1690
rect 297 -1733 330 -1690
rect 264 -1733 297 -1690
rect 363 -1733 396 -1690
rect 429 -1733 462 -1690
rect 462 -1733 495 -1690
rect 495 -1733 528 -1690
rect 561 -1733 594 -1690
rect 528 -1733 561 -1690
rect 627 -1733 660 -1690
rect 693 -1733 726 -1690
rect 660 -1733 693 -1690
rect 759 -1733 792 -1690
rect 825 -1733 858 -1690
rect 792 -1733 825 -1690
rect 891 -1733 924 -1690
rect -33 -1804 0 -1761
rect 33 -1804 66 -1761
rect 66 -1804 99 -1761
rect 99 -1804 132 -1761
rect 165 -1804 198 -1761
rect 198 -1804 231 -1761
rect 231 -1804 264 -1761
rect 297 -1804 330 -1761
rect 264 -1804 297 -1761
rect 363 -1804 396 -1761
rect 429 -1804 462 -1761
rect 396 -1804 429 -1761
rect 495 -1804 528 -1761
rect 561 -1804 594 -1761
rect 594 -1804 627 -1761
rect 627 -1804 660 -1761
rect 693 -1804 726 -1761
rect 726 -1804 759 -1761
rect 759 -1804 792 -1761
rect 825 -1804 858 -1761
rect 858 -1804 891 -1761
rect 891 -1804 924 -1761
rect -33 -1875 0 -1832
rect 33 -1875 66 -1832
rect 66 -1875 99 -1832
rect 99 -1875 132 -1832
rect 165 -1875 198 -1832
rect 198 -1875 231 -1832
rect 231 -1875 264 -1832
rect 297 -1875 330 -1832
rect 264 -1875 297 -1832
rect 363 -1875 396 -1832
rect 429 -1875 462 -1832
rect 396 -1875 429 -1832
rect 495 -1875 528 -1832
rect 561 -1875 594 -1832
rect 594 -1875 627 -1832
rect 627 -1875 660 -1832
rect 693 -1875 726 -1832
rect 726 -1875 759 -1832
rect 759 -1875 792 -1832
rect 825 -1875 858 -1832
rect 792 -1875 825 -1832
rect 891 -1875 924 -1832
rect -33 -1946 0 -1903
rect 33 -1946 66 -1903
rect 66 -1946 99 -1903
rect 99 -1946 132 -1903
rect 165 -1946 198 -1903
rect 198 -1946 231 -1903
rect 231 -1946 264 -1903
rect 297 -1946 330 -1903
rect 264 -1946 297 -1903
rect 363 -1946 396 -1903
rect 429 -1946 462 -1903
rect 396 -1946 429 -1903
rect 495 -1946 528 -1903
rect 561 -1946 594 -1903
rect 594 -1946 627 -1903
rect 627 -1946 660 -1903
rect 693 -1946 726 -1903
rect 660 -1946 693 -1903
rect 759 -1946 792 -1903
rect 825 -1946 858 -1903
rect 858 -1946 891 -1903
rect 891 -1946 924 -1903
rect -33 -2017 0 -1974
rect 33 -2017 66 -1974
rect 66 -2017 99 -1974
rect 99 -2017 132 -1974
rect 165 -2017 198 -1974
rect 198 -2017 231 -1974
rect 231 -2017 264 -1974
rect 297 -2017 330 -1974
rect 264 -2017 297 -1974
rect 363 -2017 396 -1974
rect 429 -2017 462 -1974
rect 396 -2017 429 -1974
rect 495 -2017 528 -1974
rect 561 -2017 594 -1974
rect 594 -2017 627 -1974
rect 627 -2017 660 -1974
rect 693 -2017 726 -1974
rect 660 -2017 693 -1974
rect 759 -2017 792 -1974
rect 825 -2017 858 -1974
rect 792 -2017 825 -1974
rect 891 -2017 924 -1974
rect -33 -2088 0 -2045
rect 33 -2088 66 -2045
rect 66 -2088 99 -2045
rect 99 -2088 132 -2045
rect 165 -2088 198 -2045
rect 198 -2088 231 -2045
rect 231 -2088 264 -2045
rect 297 -2088 330 -2045
rect 264 -2088 297 -2045
rect 363 -2088 396 -2045
rect 429 -2088 462 -2045
rect 396 -2088 429 -2045
rect 495 -2088 528 -2045
rect 561 -2088 594 -2045
rect 528 -2088 561 -2045
rect 627 -2088 660 -2045
rect 693 -2088 726 -2045
rect 726 -2088 759 -2045
rect 759 -2088 792 -2045
rect 825 -2088 858 -2045
rect 858 -2088 891 -2045
rect 891 -2088 924 -2045
rect -33 -2159 0 -2116
rect 33 -2159 66 -2116
rect 66 -2159 99 -2116
rect 99 -2159 132 -2116
rect 165 -2159 198 -2116
rect 198 -2159 231 -2116
rect 231 -2159 264 -2116
rect 297 -2159 330 -2116
rect 264 -2159 297 -2116
rect 363 -2159 396 -2116
rect 429 -2159 462 -2116
rect 396 -2159 429 -2116
rect 495 -2159 528 -2116
rect 561 -2159 594 -2116
rect 528 -2159 561 -2116
rect 627 -2159 660 -2116
rect 693 -2159 726 -2116
rect 726 -2159 759 -2116
rect 759 -2159 792 -2116
rect 825 -2159 858 -2116
rect 792 -2159 825 -2116
rect 891 -2159 924 -2116
rect -33 -2230 0 -2187
rect 33 -2230 66 -2187
rect 66 -2230 99 -2187
rect 99 -2230 132 -2187
rect 165 -2230 198 -2187
rect 198 -2230 231 -2187
rect 231 -2230 264 -2187
rect 297 -2230 330 -2187
rect 264 -2230 297 -2187
rect 363 -2230 396 -2187
rect 429 -2230 462 -2187
rect 396 -2230 429 -2187
rect 495 -2230 528 -2187
rect 561 -2230 594 -2187
rect 528 -2230 561 -2187
rect 627 -2230 660 -2187
rect 693 -2230 726 -2187
rect 660 -2230 693 -2187
rect 759 -2230 792 -2187
rect 825 -2230 858 -2187
rect 858 -2230 891 -2187
rect 891 -2230 924 -2187
rect -33 -2301 0 -2258
rect 33 -2301 66 -2258
rect 66 -2301 99 -2258
rect 99 -2301 132 -2258
rect 165 -2301 198 -2258
rect 198 -2301 231 -2258
rect 231 -2301 264 -2258
rect 297 -2301 330 -2258
rect 264 -2301 297 -2258
rect 363 -2301 396 -2258
rect 429 -2301 462 -2258
rect 396 -2301 429 -2258
rect 495 -2301 528 -2258
rect 561 -2301 594 -2258
rect 528 -2301 561 -2258
rect 627 -2301 660 -2258
rect 693 -2301 726 -2258
rect 660 -2301 693 -2258
rect 759 -2301 792 -2258
rect 825 -2301 858 -2258
rect 792 -2301 825 -2258
rect 891 -2301 924 -2258
rect -33 -2372 0 -2329
rect 33 -2372 66 -2329
rect 66 -2372 99 -2329
rect 99 -2372 132 -2329
rect 165 -2372 198 -2329
rect 132 -2372 165 -2329
rect 231 -2372 264 -2329
rect 297 -2372 330 -2329
rect 330 -2372 363 -2329
rect 363 -2372 396 -2329
rect 429 -2372 462 -2329
rect 462 -2372 495 -2329
rect 495 -2372 528 -2329
rect 561 -2372 594 -2329
rect 594 -2372 627 -2329
rect 627 -2372 660 -2329
rect 693 -2372 726 -2329
rect 726 -2372 759 -2329
rect 759 -2372 792 -2329
rect 825 -2372 858 -2329
rect 858 -2372 891 -2329
rect 891 -2372 924 -2329
rect -33 -2443 0 -2400
rect 33 -2443 66 -2400
rect 66 -2443 99 -2400
rect 99 -2443 132 -2400
rect 165 -2443 198 -2400
rect 132 -2443 165 -2400
rect 231 -2443 264 -2400
rect 297 -2443 330 -2400
rect 330 -2443 363 -2400
rect 363 -2443 396 -2400
rect 429 -2443 462 -2400
rect 462 -2443 495 -2400
rect 495 -2443 528 -2400
rect 561 -2443 594 -2400
rect 594 -2443 627 -2400
rect 627 -2443 660 -2400
rect 693 -2443 726 -2400
rect 726 -2443 759 -2400
rect 759 -2443 792 -2400
rect 825 -2443 858 -2400
rect 792 -2443 825 -2400
rect 891 -2443 924 -2400
rect -33 -2514 0 -2471
rect 33 -2514 66 -2471
rect 66 -2514 99 -2471
rect 99 -2514 132 -2471
rect 165 -2514 198 -2471
rect 132 -2514 165 -2471
rect 231 -2514 264 -2471
rect 297 -2514 330 -2471
rect 330 -2514 363 -2471
rect 363 -2514 396 -2471
rect 429 -2514 462 -2471
rect 462 -2514 495 -2471
rect 495 -2514 528 -2471
rect 561 -2514 594 -2471
rect 594 -2514 627 -2471
rect 627 -2514 660 -2471
rect 693 -2514 726 -2471
rect 660 -2514 693 -2471
rect 759 -2514 792 -2471
rect 825 -2514 858 -2471
rect 858 -2514 891 -2471
rect 891 -2514 924 -2471
rect -33 -2585 0 -2542
rect 33 -2585 66 -2542
rect 66 -2585 99 -2542
rect 99 -2585 132 -2542
rect 165 -2585 198 -2542
rect 132 -2585 165 -2542
rect 231 -2585 264 -2542
rect 297 -2585 330 -2542
rect 330 -2585 363 -2542
rect 363 -2585 396 -2542
rect 429 -2585 462 -2542
rect 462 -2585 495 -2542
rect 495 -2585 528 -2542
rect 561 -2585 594 -2542
rect 594 -2585 627 -2542
rect 627 -2585 660 -2542
rect 693 -2585 726 -2542
rect 660 -2585 693 -2542
rect 759 -2585 792 -2542
rect 825 -2585 858 -2542
rect 792 -2585 825 -2542
rect 891 -2585 924 -2542
rect -33 -2656 0 -2613
rect 33 -2656 66 -2613
rect 66 -2656 99 -2613
rect 99 -2656 132 -2613
rect 165 -2656 198 -2613
rect 132 -2656 165 -2613
rect 231 -2656 264 -2613
rect 297 -2656 330 -2613
rect 330 -2656 363 -2613
rect 363 -2656 396 -2613
rect 429 -2656 462 -2613
rect 462 -2656 495 -2613
rect 495 -2656 528 -2613
rect 561 -2656 594 -2613
rect 528 -2656 561 -2613
rect 627 -2656 660 -2613
rect 693 -2656 726 -2613
rect 726 -2656 759 -2613
rect 759 -2656 792 -2613
rect 825 -2656 858 -2613
rect 858 -2656 891 -2613
rect 891 -2656 924 -2613
rect -33 -2727 0 -2684
rect 33 -2727 66 -2684
rect 66 -2727 99 -2684
rect 99 -2727 132 -2684
rect 165 -2727 198 -2684
rect 132 -2727 165 -2684
rect 231 -2727 264 -2684
rect 297 -2727 330 -2684
rect 330 -2727 363 -2684
rect 363 -2727 396 -2684
rect 429 -2727 462 -2684
rect 462 -2727 495 -2684
rect 495 -2727 528 -2684
rect 561 -2727 594 -2684
rect 528 -2727 561 -2684
rect 627 -2727 660 -2684
rect 693 -2727 726 -2684
rect 726 -2727 759 -2684
rect 759 -2727 792 -2684
rect 825 -2727 858 -2684
rect 792 -2727 825 -2684
rect 891 -2727 924 -2684
rect -33 -2798 0 -2755
rect 33 -2798 66 -2755
rect 66 -2798 99 -2755
rect 99 -2798 132 -2755
rect 165 -2798 198 -2755
rect 132 -2798 165 -2755
rect 231 -2798 264 -2755
rect 297 -2798 330 -2755
rect 330 -2798 363 -2755
rect 363 -2798 396 -2755
rect 429 -2798 462 -2755
rect 462 -2798 495 -2755
rect 495 -2798 528 -2755
rect 561 -2798 594 -2755
rect 528 -2798 561 -2755
rect 627 -2798 660 -2755
rect 693 -2798 726 -2755
rect 660 -2798 693 -2755
rect 759 -2798 792 -2755
rect 825 -2798 858 -2755
rect 858 -2798 891 -2755
rect 891 -2798 924 -2755
rect -33 -2869 0 -2826
rect 33 -2869 66 -2826
rect 66 -2869 99 -2826
rect 99 -2869 132 -2826
rect 165 -2869 198 -2826
rect 132 -2869 165 -2826
rect 231 -2869 264 -2826
rect 297 -2869 330 -2826
rect 330 -2869 363 -2826
rect 363 -2869 396 -2826
rect 429 -2869 462 -2826
rect 462 -2869 495 -2826
rect 495 -2869 528 -2826
rect 561 -2869 594 -2826
rect 528 -2869 561 -2826
rect 627 -2869 660 -2826
rect 693 -2869 726 -2826
rect 660 -2869 693 -2826
rect 759 -2869 792 -2826
rect 825 -2869 858 -2826
rect 792 -2869 825 -2826
rect 891 -2869 924 -2826
rect -33 -2940 0 -2897
rect 33 -2940 66 -2897
rect 66 -2940 99 -2897
rect 99 -2940 132 -2897
rect 165 -2940 198 -2897
rect 132 -2940 165 -2897
rect 231 -2940 264 -2897
rect 297 -2940 330 -2897
rect 330 -2940 363 -2897
rect 363 -2940 396 -2897
rect 429 -2940 462 -2897
rect 396 -2940 429 -2897
rect 495 -2940 528 -2897
rect 561 -2940 594 -2897
rect 594 -2940 627 -2897
rect 627 -2940 660 -2897
rect 693 -2940 726 -2897
rect 726 -2940 759 -2897
rect 759 -2940 792 -2897
rect 825 -2940 858 -2897
rect 858 -2940 891 -2897
rect 891 -2940 924 -2897
rect -33 -3011 0 -2968
rect 33 -3011 66 -2968
rect 66 -3011 99 -2968
rect 99 -3011 132 -2968
rect 165 -3011 198 -2968
rect 132 -3011 165 -2968
rect 231 -3011 264 -2968
rect 297 -3011 330 -2968
rect 330 -3011 363 -2968
rect 363 -3011 396 -2968
rect 429 -3011 462 -2968
rect 396 -3011 429 -2968
rect 495 -3011 528 -2968
rect 561 -3011 594 -2968
rect 594 -3011 627 -2968
rect 627 -3011 660 -2968
rect 693 -3011 726 -2968
rect 726 -3011 759 -2968
rect 759 -3011 792 -2968
rect 825 -3011 858 -2968
rect 792 -3011 825 -2968
rect 891 -3011 924 -2968
rect -33 -3082 0 -3039
rect 33 -3082 66 -3039
rect 66 -3082 99 -3039
rect 99 -3082 132 -3039
rect 165 -3082 198 -3039
rect 132 -3082 165 -3039
rect 231 -3082 264 -3039
rect 297 -3082 330 -3039
rect 330 -3082 363 -3039
rect 363 -3082 396 -3039
rect 429 -3082 462 -3039
rect 396 -3082 429 -3039
rect 495 -3082 528 -3039
rect 561 -3082 594 -3039
rect 594 -3082 627 -3039
rect 627 -3082 660 -3039
rect 693 -3082 726 -3039
rect 660 -3082 693 -3039
rect 759 -3082 792 -3039
rect 825 -3082 858 -3039
rect 858 -3082 891 -3039
rect 891 -3082 924 -3039
rect -33 -3153 0 -3110
rect 33 -3153 66 -3110
rect 66 -3153 99 -3110
rect 99 -3153 132 -3110
rect 165 -3153 198 -3110
rect 132 -3153 165 -3110
rect 231 -3153 264 -3110
rect 297 -3153 330 -3110
rect 330 -3153 363 -3110
rect 363 -3153 396 -3110
rect 429 -3153 462 -3110
rect 396 -3153 429 -3110
rect 495 -3153 528 -3110
rect 561 -3153 594 -3110
rect 594 -3153 627 -3110
rect 627 -3153 660 -3110
rect 693 -3153 726 -3110
rect 660 -3153 693 -3110
rect 759 -3153 792 -3110
rect 825 -3153 858 -3110
rect 792 -3153 825 -3110
rect 891 -3153 924 -3110
rect -33 -3224 0 -3181
rect 33 -3224 66 -3181
rect 66 -3224 99 -3181
rect 99 -3224 132 -3181
rect 165 -3224 198 -3181
rect 132 -3224 165 -3181
rect 231 -3224 264 -3181
rect 297 -3224 330 -3181
rect 330 -3224 363 -3181
rect 363 -3224 396 -3181
rect 429 -3224 462 -3181
rect 396 -3224 429 -3181
rect 495 -3224 528 -3181
rect 561 -3224 594 -3181
rect 528 -3224 561 -3181
rect 627 -3224 660 -3181
rect 693 -3224 726 -3181
rect 726 -3224 759 -3181
rect 759 -3224 792 -3181
rect 825 -3224 858 -3181
rect 858 -3224 891 -3181
rect 891 -3224 924 -3181
rect -33 -3295 0 -3252
rect 33 -3295 66 -3252
rect 66 -3295 99 -3252
rect 99 -3295 132 -3252
rect 165 -3295 198 -3252
rect 132 -3295 165 -3252
rect 231 -3295 264 -3252
rect 297 -3295 330 -3252
rect 330 -3295 363 -3252
rect 363 -3295 396 -3252
rect 429 -3295 462 -3252
rect 396 -3295 429 -3252
rect 495 -3295 528 -3252
rect 561 -3295 594 -3252
rect 528 -3295 561 -3252
rect 627 -3295 660 -3252
rect 693 -3295 726 -3252
rect 726 -3295 759 -3252
rect 759 -3295 792 -3252
rect 825 -3295 858 -3252
rect 792 -3295 825 -3252
rect 891 -3295 924 -3252
rect -33 -3366 0 -3323
rect 33 -3366 66 -3323
rect 66 -3366 99 -3323
rect 99 -3366 132 -3323
rect 165 -3366 198 -3323
rect 132 -3366 165 -3323
rect 231 -3366 264 -3323
rect 297 -3366 330 -3323
rect 330 -3366 363 -3323
rect 363 -3366 396 -3323
rect 429 -3366 462 -3323
rect 396 -3366 429 -3323
rect 495 -3366 528 -3323
rect 561 -3366 594 -3323
rect 528 -3366 561 -3323
rect 627 -3366 660 -3323
rect 693 -3366 726 -3323
rect 660 -3366 693 -3323
rect 759 -3366 792 -3323
rect 825 -3366 858 -3323
rect 858 -3366 891 -3323
rect 891 -3366 924 -3323
rect -33 -3437 0 -3394
rect 33 -3437 66 -3394
rect 66 -3437 99 -3394
rect 99 -3437 132 -3394
rect 165 -3437 198 -3394
rect 132 -3437 165 -3394
rect 231 -3437 264 -3394
rect 297 -3437 330 -3394
rect 330 -3437 363 -3394
rect 363 -3437 396 -3394
rect 429 -3437 462 -3394
rect 396 -3437 429 -3394
rect 495 -3437 528 -3394
rect 561 -3437 594 -3394
rect 528 -3437 561 -3394
rect 627 -3437 660 -3394
rect 693 -3437 726 -3394
rect 660 -3437 693 -3394
rect 759 -3437 792 -3394
rect 825 -3437 858 -3394
rect 792 -3437 825 -3394
rect 891 -3437 924 -3394
rect -33 -3508 0 -3465
rect 33 -3508 66 -3465
rect 66 -3508 99 -3465
rect 99 -3508 132 -3465
rect 165 -3508 198 -3465
rect 132 -3508 165 -3465
rect 231 -3508 264 -3465
rect 297 -3508 330 -3465
rect 264 -3508 297 -3465
rect 363 -3508 396 -3465
rect 429 -3508 462 -3465
rect 462 -3508 495 -3465
rect 495 -3508 528 -3465
rect 561 -3508 594 -3465
rect 594 -3508 627 -3465
rect 627 -3508 660 -3465
rect 693 -3508 726 -3465
rect 726 -3508 759 -3465
rect 759 -3508 792 -3465
rect 825 -3508 858 -3465
rect 858 -3508 891 -3465
rect 891 -3508 924 -3465
rect -33 -3579 0 -3536
rect 33 -3579 66 -3536
rect 66 -3579 99 -3536
rect 99 -3579 132 -3536
rect 165 -3579 198 -3536
rect 132 -3579 165 -3536
rect 231 -3579 264 -3536
rect 297 -3579 330 -3536
rect 264 -3579 297 -3536
rect 363 -3579 396 -3536
rect 429 -3579 462 -3536
rect 462 -3579 495 -3536
rect 495 -3579 528 -3536
rect 561 -3579 594 -3536
rect 594 -3579 627 -3536
rect 627 -3579 660 -3536
rect 693 -3579 726 -3536
rect 726 -3579 759 -3536
rect 759 -3579 792 -3536
rect 825 -3579 858 -3536
rect 792 -3579 825 -3536
rect 891 -3579 924 -3536
rect -33 -3650 0 -3607
rect 33 -3650 66 -3607
rect 66 -3650 99 -3607
rect 99 -3650 132 -3607
rect 165 -3650 198 -3607
rect 132 -3650 165 -3607
rect 231 -3650 264 -3607
rect 297 -3650 330 -3607
rect 264 -3650 297 -3607
rect 363 -3650 396 -3607
rect 429 -3650 462 -3607
rect 462 -3650 495 -3607
rect 495 -3650 528 -3607
rect 561 -3650 594 -3607
rect 594 -3650 627 -3607
rect 627 -3650 660 -3607
rect 693 -3650 726 -3607
rect 660 -3650 693 -3607
rect 759 -3650 792 -3607
rect 825 -3650 858 -3607
rect 858 -3650 891 -3607
rect 891 -3650 924 -3607
rect -33 -3721 0 -3678
rect 33 -3721 66 -3678
rect 66 -3721 99 -3678
rect 99 -3721 132 -3678
rect 165 -3721 198 -3678
rect 132 -3721 165 -3678
rect 231 -3721 264 -3678
rect 297 -3721 330 -3678
rect 264 -3721 297 -3678
rect 363 -3721 396 -3678
rect 429 -3721 462 -3678
rect 462 -3721 495 -3678
rect 495 -3721 528 -3678
rect 561 -3721 594 -3678
rect 594 -3721 627 -3678
rect 627 -3721 660 -3678
rect 693 -3721 726 -3678
rect 660 -3721 693 -3678
rect 759 -3721 792 -3678
rect 825 -3721 858 -3678
rect 792 -3721 825 -3678
rect 891 -3721 924 -3678
rect -33 -3792 0 -3749
rect 33 -3792 66 -3749
rect 66 -3792 99 -3749
rect 99 -3792 132 -3749
rect 165 -3792 198 -3749
rect 132 -3792 165 -3749
rect 231 -3792 264 -3749
rect 297 -3792 330 -3749
rect 264 -3792 297 -3749
rect 363 -3792 396 -3749
rect 429 -3792 462 -3749
rect 462 -3792 495 -3749
rect 495 -3792 528 -3749
rect 561 -3792 594 -3749
rect 528 -3792 561 -3749
rect 627 -3792 660 -3749
rect 693 -3792 726 -3749
rect 726 -3792 759 -3749
rect 759 -3792 792 -3749
rect 825 -3792 858 -3749
rect 858 -3792 891 -3749
rect 891 -3792 924 -3749
rect -33 -3863 0 -3820
rect 33 -3863 66 -3820
rect 66 -3863 99 -3820
rect 99 -3863 132 -3820
rect 165 -3863 198 -3820
rect 132 -3863 165 -3820
rect 231 -3863 264 -3820
rect 297 -3863 330 -3820
rect 264 -3863 297 -3820
rect 363 -3863 396 -3820
rect 429 -3863 462 -3820
rect 462 -3863 495 -3820
rect 495 -3863 528 -3820
rect 561 -3863 594 -3820
rect 528 -3863 561 -3820
rect 627 -3863 660 -3820
rect 693 -3863 726 -3820
rect 726 -3863 759 -3820
rect 759 -3863 792 -3820
rect 825 -3863 858 -3820
rect 792 -3863 825 -3820
rect 891 -3863 924 -3820
rect -33 -3934 0 -3891
rect 33 -3934 66 -3891
rect 66 -3934 99 -3891
rect 99 -3934 132 -3891
rect 165 -3934 198 -3891
rect 132 -3934 165 -3891
rect 231 -3934 264 -3891
rect 297 -3934 330 -3891
rect 264 -3934 297 -3891
rect 363 -3934 396 -3891
rect 429 -3934 462 -3891
rect 462 -3934 495 -3891
rect 495 -3934 528 -3891
rect 561 -3934 594 -3891
rect 528 -3934 561 -3891
rect 627 -3934 660 -3891
rect 693 -3934 726 -3891
rect 660 -3934 693 -3891
rect 759 -3934 792 -3891
rect 825 -3934 858 -3891
rect 858 -3934 891 -3891
rect 891 -3934 924 -3891
rect -33 -4005 0 -3962
rect 33 -4005 66 -3962
rect 66 -4005 99 -3962
rect 99 -4005 132 -3962
rect 165 -4005 198 -3962
rect 132 -4005 165 -3962
rect 231 -4005 264 -3962
rect 297 -4005 330 -3962
rect 264 -4005 297 -3962
rect 363 -4005 396 -3962
rect 429 -4005 462 -3962
rect 462 -4005 495 -3962
rect 495 -4005 528 -3962
rect 561 -4005 594 -3962
rect 528 -4005 561 -3962
rect 627 -4005 660 -3962
rect 693 -4005 726 -3962
rect 660 -4005 693 -3962
rect 759 -4005 792 -3962
rect 825 -4005 858 -3962
rect 792 -4005 825 -3962
rect 891 -4005 924 -3962
rect -33 -4076 0 -4033
rect 33 -4076 66 -4033
rect 66 -4076 99 -4033
rect 99 -4076 132 -4033
rect 165 -4076 198 -4033
rect 132 -4076 165 -4033
rect 231 -4076 264 -4033
rect 297 -4076 330 -4033
rect 264 -4076 297 -4033
rect 363 -4076 396 -4033
rect 429 -4076 462 -4033
rect 396 -4076 429 -4033
rect 495 -4076 528 -4033
rect 561 -4076 594 -4033
rect 594 -4076 627 -4033
rect 627 -4076 660 -4033
rect 693 -4076 726 -4033
rect 726 -4076 759 -4033
rect 759 -4076 792 -4033
rect 825 -4076 858 -4033
rect 858 -4076 891 -4033
rect 891 -4076 924 -4033
rect -33 -4147 0 -4104
rect 33 -4147 66 -4104
rect 66 -4147 99 -4104
rect 99 -4147 132 -4104
rect 165 -4147 198 -4104
rect 132 -4147 165 -4104
rect 231 -4147 264 -4104
rect 297 -4147 330 -4104
rect 264 -4147 297 -4104
rect 363 -4147 396 -4104
rect 429 -4147 462 -4104
rect 396 -4147 429 -4104
rect 495 -4147 528 -4104
rect 561 -4147 594 -4104
rect 594 -4147 627 -4104
rect 627 -4147 660 -4104
rect 693 -4147 726 -4104
rect 726 -4147 759 -4104
rect 759 -4147 792 -4104
rect 825 -4147 858 -4104
rect 792 -4147 825 -4104
rect 891 -4147 924 -4104
rect -33 -4218 0 -4175
rect 33 -4218 66 -4175
rect 66 -4218 99 -4175
rect 99 -4218 132 -4175
rect 165 -4218 198 -4175
rect 132 -4218 165 -4175
rect 231 -4218 264 -4175
rect 297 -4218 330 -4175
rect 264 -4218 297 -4175
rect 363 -4218 396 -4175
rect 429 -4218 462 -4175
rect 396 -4218 429 -4175
rect 495 -4218 528 -4175
rect 561 -4218 594 -4175
rect 594 -4218 627 -4175
rect 627 -4218 660 -4175
rect 693 -4218 726 -4175
rect 660 -4218 693 -4175
rect 759 -4218 792 -4175
rect 825 -4218 858 -4175
rect 858 -4218 891 -4175
rect 891 -4218 924 -4175
rect -33 -4289 0 -4246
rect 33 -4289 66 -4246
rect 66 -4289 99 -4246
rect 99 -4289 132 -4246
rect 165 -4289 198 -4246
rect 132 -4289 165 -4246
rect 231 -4289 264 -4246
rect 297 -4289 330 -4246
rect 264 -4289 297 -4246
rect 363 -4289 396 -4246
rect 429 -4289 462 -4246
rect 396 -4289 429 -4246
rect 495 -4289 528 -4246
rect 561 -4289 594 -4246
rect 594 -4289 627 -4246
rect 627 -4289 660 -4246
rect 693 -4289 726 -4246
rect 660 -4289 693 -4246
rect 759 -4289 792 -4246
rect 825 -4289 858 -4246
rect 792 -4289 825 -4246
rect 891 -4289 924 -4246
rect -33 -4360 0 -4317
rect 33 -4360 66 -4317
rect 66 -4360 99 -4317
rect 99 -4360 132 -4317
rect 165 -4360 198 -4317
rect 132 -4360 165 -4317
rect 231 -4360 264 -4317
rect 297 -4360 330 -4317
rect 264 -4360 297 -4317
rect 363 -4360 396 -4317
rect 429 -4360 462 -4317
rect 396 -4360 429 -4317
rect 495 -4360 528 -4317
rect 561 -4360 594 -4317
rect 528 -4360 561 -4317
rect 627 -4360 660 -4317
rect 693 -4360 726 -4317
rect 726 -4360 759 -4317
rect 759 -4360 792 -4317
rect 825 -4360 858 -4317
rect 858 -4360 891 -4317
rect 891 -4360 924 -4317
rect -33 -4431 0 -4388
rect 33 -4431 66 -4388
rect 66 -4431 99 -4388
rect 99 -4431 132 -4388
rect 165 -4431 198 -4388
rect 132 -4431 165 -4388
rect 231 -4431 264 -4388
rect 297 -4431 330 -4388
rect 264 -4431 297 -4388
rect 363 -4431 396 -4388
rect 429 -4431 462 -4388
rect 396 -4431 429 -4388
rect 495 -4431 528 -4388
rect 561 -4431 594 -4388
rect 528 -4431 561 -4388
rect 627 -4431 660 -4388
rect 693 -4431 726 -4388
rect 726 -4431 759 -4388
rect 759 -4431 792 -4388
rect 825 -4431 858 -4388
rect 792 -4431 825 -4388
rect 891 -4431 924 -4388
rect -33 -4502 0 -4459
rect 33 -4502 66 -4459
rect 66 -4502 99 -4459
rect 99 -4502 132 -4459
rect 165 -4502 198 -4459
rect 132 -4502 165 -4459
rect 231 -4502 264 -4459
rect 297 -4502 330 -4459
rect 264 -4502 297 -4459
rect 363 -4502 396 -4459
rect 429 -4502 462 -4459
rect 396 -4502 429 -4459
rect 495 -4502 528 -4459
rect 561 -4502 594 -4459
rect 528 -4502 561 -4459
rect 627 -4502 660 -4459
rect 693 -4502 726 -4459
rect 660 -4502 693 -4459
rect 759 -4502 792 -4459
rect 825 -4502 858 -4459
rect 858 -4502 891 -4459
rect 891 -4502 924 -4459
rect -33 -4573 0 -4530
rect 33 -4573 66 -4530
rect 66 -4573 99 -4530
rect 99 -4573 132 -4530
rect 165 -4573 198 -4530
rect 132 -4573 165 -4530
rect 231 -4573 264 -4530
rect 297 -4573 330 -4530
rect 264 -4573 297 -4530
rect 363 -4573 396 -4530
rect 429 -4573 462 -4530
rect 396 -4573 429 -4530
rect 495 -4573 528 -4530
rect 561 -4573 594 -4530
rect 528 -4573 561 -4530
rect 627 -4573 660 -4530
rect 693 -4573 726 -4530
rect 660 -4573 693 -4530
rect 759 -4573 792 -4530
rect 825 -4573 858 -4530
rect 792 -4573 825 -4530
rect 891 -4573 924 -4530
rect -33 -4644 0 -4601
rect 33 -4644 66 -4601
rect 0 -4644 33 -4601
rect 99 -4644 132 -4601
rect 165 -4644 198 -4601
rect 198 -4644 231 -4601
rect 231 -4644 264 -4601
rect 297 -4644 330 -4601
rect 330 -4644 363 -4601
rect 363 -4644 396 -4601
rect 429 -4644 462 -4601
rect 462 -4644 495 -4601
rect 495 -4644 528 -4601
rect 561 -4644 594 -4601
rect 594 -4644 627 -4601
rect 627 -4644 660 -4601
rect 693 -4644 726 -4601
rect 726 -4644 759 -4601
rect 759 -4644 792 -4601
rect 825 -4644 858 -4601
rect 858 -4644 891 -4601
rect 891 -4644 924 -4601
rect -33 -4715 0 -4672
rect 33 -4715 66 -4672
rect 0 -4715 33 -4672
rect 99 -4715 132 -4672
rect 165 -4715 198 -4672
rect 198 -4715 231 -4672
rect 231 -4715 264 -4672
rect 297 -4715 330 -4672
rect 330 -4715 363 -4672
rect 363 -4715 396 -4672
rect 429 -4715 462 -4672
rect 462 -4715 495 -4672
rect 495 -4715 528 -4672
rect 561 -4715 594 -4672
rect 594 -4715 627 -4672
rect 627 -4715 660 -4672
rect 693 -4715 726 -4672
rect 726 -4715 759 -4672
rect 759 -4715 792 -4672
rect 825 -4715 858 -4672
rect 792 -4715 825 -4672
rect 891 -4715 924 -4672
rect -33 -4786 0 -4743
rect 33 -4786 66 -4743
rect 0 -4786 33 -4743
rect 99 -4786 132 -4743
rect 165 -4786 198 -4743
rect 198 -4786 231 -4743
rect 231 -4786 264 -4743
rect 297 -4786 330 -4743
rect 330 -4786 363 -4743
rect 363 -4786 396 -4743
rect 429 -4786 462 -4743
rect 462 -4786 495 -4743
rect 495 -4786 528 -4743
rect 561 -4786 594 -4743
rect 594 -4786 627 -4743
rect 627 -4786 660 -4743
rect 693 -4786 726 -4743
rect 660 -4786 693 -4743
rect 759 -4786 792 -4743
rect 825 -4786 858 -4743
rect 858 -4786 891 -4743
rect 891 -4786 924 -4743
rect -33 -4857 0 -4814
rect 33 -4857 66 -4814
rect 0 -4857 33 -4814
rect 99 -4857 132 -4814
rect 165 -4857 198 -4814
rect 198 -4857 231 -4814
rect 231 -4857 264 -4814
rect 297 -4857 330 -4814
rect 330 -4857 363 -4814
rect 363 -4857 396 -4814
rect 429 -4857 462 -4814
rect 462 -4857 495 -4814
rect 495 -4857 528 -4814
rect 561 -4857 594 -4814
rect 594 -4857 627 -4814
rect 627 -4857 660 -4814
rect 693 -4857 726 -4814
rect 660 -4857 693 -4814
rect 759 -4857 792 -4814
rect 825 -4857 858 -4814
rect 792 -4857 825 -4814
rect 891 -4857 924 -4814
rect -33 -4928 0 -4885
rect 33 -4928 66 -4885
rect 0 -4928 33 -4885
rect 99 -4928 132 -4885
rect 165 -4928 198 -4885
rect 198 -4928 231 -4885
rect 231 -4928 264 -4885
rect 297 -4928 330 -4885
rect 330 -4928 363 -4885
rect 363 -4928 396 -4885
rect 429 -4928 462 -4885
rect 462 -4928 495 -4885
rect 495 -4928 528 -4885
rect 561 -4928 594 -4885
rect 528 -4928 561 -4885
rect 627 -4928 660 -4885
rect 693 -4928 726 -4885
rect 726 -4928 759 -4885
rect 759 -4928 792 -4885
rect 825 -4928 858 -4885
rect 858 -4928 891 -4885
rect 891 -4928 924 -4885
rect -33 -4999 0 -4956
rect 33 -4999 66 -4956
rect 0 -4999 33 -4956
rect 99 -4999 132 -4956
rect 165 -4999 198 -4956
rect 198 -4999 231 -4956
rect 231 -4999 264 -4956
rect 297 -4999 330 -4956
rect 330 -4999 363 -4956
rect 363 -4999 396 -4956
rect 429 -4999 462 -4956
rect 462 -4999 495 -4956
rect 495 -4999 528 -4956
rect 561 -4999 594 -4956
rect 528 -4999 561 -4956
rect 627 -4999 660 -4956
rect 693 -4999 726 -4956
rect 726 -4999 759 -4956
rect 759 -4999 792 -4956
rect 825 -4999 858 -4956
rect 792 -4999 825 -4956
rect 891 -4999 924 -4956
rect -33 -5070 0 -5027
rect 33 -5070 66 -5027
rect 0 -5070 33 -5027
rect 99 -5070 132 -5027
rect 165 -5070 198 -5027
rect 198 -5070 231 -5027
rect 231 -5070 264 -5027
rect 297 -5070 330 -5027
rect 330 -5070 363 -5027
rect 363 -5070 396 -5027
rect 429 -5070 462 -5027
rect 462 -5070 495 -5027
rect 495 -5070 528 -5027
rect 561 -5070 594 -5027
rect 528 -5070 561 -5027
rect 627 -5070 660 -5027
rect 693 -5070 726 -5027
rect 660 -5070 693 -5027
rect 759 -5070 792 -5027
rect 825 -5070 858 -5027
rect 858 -5070 891 -5027
rect 891 -5070 924 -5027
rect -33 -5141 0 -5098
rect 33 -5141 66 -5098
rect 0 -5141 33 -5098
rect 99 -5141 132 -5098
rect 165 -5141 198 -5098
rect 198 -5141 231 -5098
rect 231 -5141 264 -5098
rect 297 -5141 330 -5098
rect 330 -5141 363 -5098
rect 363 -5141 396 -5098
rect 429 -5141 462 -5098
rect 462 -5141 495 -5098
rect 495 -5141 528 -5098
rect 561 -5141 594 -5098
rect 528 -5141 561 -5098
rect 627 -5141 660 -5098
rect 693 -5141 726 -5098
rect 660 -5141 693 -5098
rect 759 -5141 792 -5098
rect 825 -5141 858 -5098
rect 792 -5141 825 -5098
rect 891 -5141 924 -5098
rect -33 -5212 0 -5169
rect 33 -5212 66 -5169
rect 0 -5212 33 -5169
rect 99 -5212 132 -5169
rect 165 -5212 198 -5169
rect 198 -5212 231 -5169
rect 231 -5212 264 -5169
rect 297 -5212 330 -5169
rect 330 -5212 363 -5169
rect 363 -5212 396 -5169
rect 429 -5212 462 -5169
rect 396 -5212 429 -5169
rect 495 -5212 528 -5169
rect 561 -5212 594 -5169
rect 594 -5212 627 -5169
rect 627 -5212 660 -5169
rect 693 -5212 726 -5169
rect 726 -5212 759 -5169
rect 759 -5212 792 -5169
rect 825 -5212 858 -5169
rect 858 -5212 891 -5169
rect 891 -5212 924 -5169
rect -33 -5283 0 -5240
rect 33 -5283 66 -5240
rect 0 -5283 33 -5240
rect 99 -5283 132 -5240
rect 165 -5283 198 -5240
rect 198 -5283 231 -5240
rect 231 -5283 264 -5240
rect 297 -5283 330 -5240
rect 330 -5283 363 -5240
rect 363 -5283 396 -5240
rect 429 -5283 462 -5240
rect 396 -5283 429 -5240
rect 495 -5283 528 -5240
rect 561 -5283 594 -5240
rect 594 -5283 627 -5240
rect 627 -5283 660 -5240
rect 693 -5283 726 -5240
rect 726 -5283 759 -5240
rect 759 -5283 792 -5240
rect 825 -5283 858 -5240
rect 792 -5283 825 -5240
rect 891 -5283 924 -5240
rect -33 -5354 0 -5311
rect 33 -5354 66 -5311
rect 0 -5354 33 -5311
rect 99 -5354 132 -5311
rect 165 -5354 198 -5311
rect 198 -5354 231 -5311
rect 231 -5354 264 -5311
rect 297 -5354 330 -5311
rect 330 -5354 363 -5311
rect 363 -5354 396 -5311
rect 429 -5354 462 -5311
rect 396 -5354 429 -5311
rect 495 -5354 528 -5311
rect 561 -5354 594 -5311
rect 594 -5354 627 -5311
rect 627 -5354 660 -5311
rect 693 -5354 726 -5311
rect 660 -5354 693 -5311
rect 759 -5354 792 -5311
rect 825 -5354 858 -5311
rect 858 -5354 891 -5311
rect 891 -5354 924 -5311
rect -33 -5425 0 -5382
rect 33 -5425 66 -5382
rect 0 -5425 33 -5382
rect 99 -5425 132 -5382
rect 165 -5425 198 -5382
rect 198 -5425 231 -5382
rect 231 -5425 264 -5382
rect 297 -5425 330 -5382
rect 330 -5425 363 -5382
rect 363 -5425 396 -5382
rect 429 -5425 462 -5382
rect 396 -5425 429 -5382
rect 495 -5425 528 -5382
rect 561 -5425 594 -5382
rect 594 -5425 627 -5382
rect 627 -5425 660 -5382
rect 693 -5425 726 -5382
rect 660 -5425 693 -5382
rect 759 -5425 792 -5382
rect 825 -5425 858 -5382
rect 792 -5425 825 -5382
rect 891 -5425 924 -5382
rect -33 -5496 0 -5453
rect 33 -5496 66 -5453
rect 0 -5496 33 -5453
rect 99 -5496 132 -5453
rect 165 -5496 198 -5453
rect 198 -5496 231 -5453
rect 231 -5496 264 -5453
rect 297 -5496 330 -5453
rect 330 -5496 363 -5453
rect 363 -5496 396 -5453
rect 429 -5496 462 -5453
rect 396 -5496 429 -5453
rect 495 -5496 528 -5453
rect 561 -5496 594 -5453
rect 528 -5496 561 -5453
rect 627 -5496 660 -5453
rect 693 -5496 726 -5453
rect 726 -5496 759 -5453
rect 759 -5496 792 -5453
rect 825 -5496 858 -5453
rect 858 -5496 891 -5453
rect 891 -5496 924 -5453
rect -33 -5567 0 -5524
rect 33 -5567 66 -5524
rect 0 -5567 33 -5524
rect 99 -5567 132 -5524
rect 165 -5567 198 -5524
rect 198 -5567 231 -5524
rect 231 -5567 264 -5524
rect 297 -5567 330 -5524
rect 330 -5567 363 -5524
rect 363 -5567 396 -5524
rect 429 -5567 462 -5524
rect 396 -5567 429 -5524
rect 495 -5567 528 -5524
rect 561 -5567 594 -5524
rect 528 -5567 561 -5524
rect 627 -5567 660 -5524
rect 693 -5567 726 -5524
rect 726 -5567 759 -5524
rect 759 -5567 792 -5524
rect 825 -5567 858 -5524
rect 792 -5567 825 -5524
rect 891 -5567 924 -5524
rect -33 -5638 0 -5595
rect 33 -5638 66 -5595
rect 0 -5638 33 -5595
rect 99 -5638 132 -5595
rect 165 -5638 198 -5595
rect 198 -5638 231 -5595
rect 231 -5638 264 -5595
rect 297 -5638 330 -5595
rect 330 -5638 363 -5595
rect 363 -5638 396 -5595
rect 429 -5638 462 -5595
rect 396 -5638 429 -5595
rect 495 -5638 528 -5595
rect 561 -5638 594 -5595
rect 528 -5638 561 -5595
rect 627 -5638 660 -5595
rect 693 -5638 726 -5595
rect 660 -5638 693 -5595
rect 759 -5638 792 -5595
rect 825 -5638 858 -5595
rect 858 -5638 891 -5595
rect 891 -5638 924 -5595
rect -33 -5709 0 -5666
rect 33 -5709 66 -5666
rect 0 -5709 33 -5666
rect 99 -5709 132 -5666
rect 165 -5709 198 -5666
rect 198 -5709 231 -5666
rect 231 -5709 264 -5666
rect 297 -5709 330 -5666
rect 330 -5709 363 -5666
rect 363 -5709 396 -5666
rect 429 -5709 462 -5666
rect 396 -5709 429 -5666
rect 495 -5709 528 -5666
rect 561 -5709 594 -5666
rect 528 -5709 561 -5666
rect 627 -5709 660 -5666
rect 693 -5709 726 -5666
rect 660 -5709 693 -5666
rect 759 -5709 792 -5666
rect 825 -5709 858 -5666
rect 792 -5709 825 -5666
rect 891 -5709 924 -5666
rect -33 -5780 0 -5737
rect 33 -5780 66 -5737
rect 0 -5780 33 -5737
rect 99 -5780 132 -5737
rect 165 -5780 198 -5737
rect 198 -5780 231 -5737
rect 231 -5780 264 -5737
rect 297 -5780 330 -5737
rect 264 -5780 297 -5737
rect 363 -5780 396 -5737
rect 429 -5780 462 -5737
rect 462 -5780 495 -5737
rect 495 -5780 528 -5737
rect 561 -5780 594 -5737
rect 594 -5780 627 -5737
rect 627 -5780 660 -5737
rect 693 -5780 726 -5737
rect 726 -5780 759 -5737
rect 759 -5780 792 -5737
rect 825 -5780 858 -5737
rect 858 -5780 891 -5737
rect 891 -5780 924 -5737
rect -33 -5851 0 -5808
rect 33 -5851 66 -5808
rect 0 -5851 33 -5808
rect 99 -5851 132 -5808
rect 165 -5851 198 -5808
rect 198 -5851 231 -5808
rect 231 -5851 264 -5808
rect 297 -5851 330 -5808
rect 264 -5851 297 -5808
rect 363 -5851 396 -5808
rect 429 -5851 462 -5808
rect 462 -5851 495 -5808
rect 495 -5851 528 -5808
rect 561 -5851 594 -5808
rect 594 -5851 627 -5808
rect 627 -5851 660 -5808
rect 693 -5851 726 -5808
rect 726 -5851 759 -5808
rect 759 -5851 792 -5808
rect 825 -5851 858 -5808
rect 792 -5851 825 -5808
rect 891 -5851 924 -5808
rect -33 -5922 0 -5879
rect 33 -5922 66 -5879
rect 0 -5922 33 -5879
rect 99 -5922 132 -5879
rect 165 -5922 198 -5879
rect 198 -5922 231 -5879
rect 231 -5922 264 -5879
rect 297 -5922 330 -5879
rect 264 -5922 297 -5879
rect 363 -5922 396 -5879
rect 429 -5922 462 -5879
rect 462 -5922 495 -5879
rect 495 -5922 528 -5879
rect 561 -5922 594 -5879
rect 594 -5922 627 -5879
rect 627 -5922 660 -5879
rect 693 -5922 726 -5879
rect 660 -5922 693 -5879
rect 759 -5922 792 -5879
rect 825 -5922 858 -5879
rect 858 -5922 891 -5879
rect 891 -5922 924 -5879
rect -33 -5993 0 -5950
rect 33 -5993 66 -5950
rect 0 -5993 33 -5950
rect 99 -5993 132 -5950
rect 165 -5993 198 -5950
rect 198 -5993 231 -5950
rect 231 -5993 264 -5950
rect 297 -5993 330 -5950
rect 264 -5993 297 -5950
rect 363 -5993 396 -5950
rect 429 -5993 462 -5950
rect 462 -5993 495 -5950
rect 495 -5993 528 -5950
rect 561 -5993 594 -5950
rect 594 -5993 627 -5950
rect 627 -5993 660 -5950
rect 693 -5993 726 -5950
rect 660 -5993 693 -5950
rect 759 -5993 792 -5950
rect 825 -5993 858 -5950
rect 792 -5993 825 -5950
rect 891 -5993 924 -5950
rect -33 -6064 0 -6021
rect 33 -6064 66 -6021
rect 0 -6064 33 -6021
rect 99 -6064 132 -6021
rect 165 -6064 198 -6021
rect 198 -6064 231 -6021
rect 231 -6064 264 -6021
rect 297 -6064 330 -6021
rect 264 -6064 297 -6021
rect 363 -6064 396 -6021
rect 429 -6064 462 -6021
rect 462 -6064 495 -6021
rect 495 -6064 528 -6021
rect 561 -6064 594 -6021
rect 528 -6064 561 -6021
rect 627 -6064 660 -6021
rect 693 -6064 726 -6021
rect 726 -6064 759 -6021
rect 759 -6064 792 -6021
rect 825 -6064 858 -6021
rect 858 -6064 891 -6021
rect 891 -6064 924 -6021
rect -33 -6135 0 -6092
rect 33 -6135 66 -6092
rect 0 -6135 33 -6092
rect 99 -6135 132 -6092
rect 165 -6135 198 -6092
rect 198 -6135 231 -6092
rect 231 -6135 264 -6092
rect 297 -6135 330 -6092
rect 264 -6135 297 -6092
rect 363 -6135 396 -6092
rect 429 -6135 462 -6092
rect 462 -6135 495 -6092
rect 495 -6135 528 -6092
rect 561 -6135 594 -6092
rect 528 -6135 561 -6092
rect 627 -6135 660 -6092
rect 693 -6135 726 -6092
rect 726 -6135 759 -6092
rect 759 -6135 792 -6092
rect 825 -6135 858 -6092
rect 792 -6135 825 -6092
rect 891 -6135 924 -6092
rect -33 -6206 0 -6163
rect 33 -6206 66 -6163
rect 0 -6206 33 -6163
rect 99 -6206 132 -6163
rect 165 -6206 198 -6163
rect 198 -6206 231 -6163
rect 231 -6206 264 -6163
rect 297 -6206 330 -6163
rect 264 -6206 297 -6163
rect 363 -6206 396 -6163
rect 429 -6206 462 -6163
rect 462 -6206 495 -6163
rect 495 -6206 528 -6163
rect 561 -6206 594 -6163
rect 528 -6206 561 -6163
rect 627 -6206 660 -6163
rect 693 -6206 726 -6163
rect 660 -6206 693 -6163
rect 759 -6206 792 -6163
rect 825 -6206 858 -6163
rect 858 -6206 891 -6163
rect 891 -6206 924 -6163
rect -33 -6277 0 -6234
rect 33 -6277 66 -6234
rect 0 -6277 33 -6234
rect 99 -6277 132 -6234
rect 165 -6277 198 -6234
rect 198 -6277 231 -6234
rect 231 -6277 264 -6234
rect 297 -6277 330 -6234
rect 264 -6277 297 -6234
rect 363 -6277 396 -6234
rect 429 -6277 462 -6234
rect 462 -6277 495 -6234
rect 495 -6277 528 -6234
rect 561 -6277 594 -6234
rect 528 -6277 561 -6234
rect 627 -6277 660 -6234
rect 693 -6277 726 -6234
rect 660 -6277 693 -6234
rect 759 -6277 792 -6234
rect 825 -6277 858 -6234
rect 792 -6277 825 -6234
rect 891 -6277 924 -6234
rect -33 -6348 0 -6305
rect 33 -6348 66 -6305
rect 0 -6348 33 -6305
rect 99 -6348 132 -6305
rect 165 -6348 198 -6305
rect 198 -6348 231 -6305
rect 231 -6348 264 -6305
rect 297 -6348 330 -6305
rect 264 -6348 297 -6305
rect 363 -6348 396 -6305
rect 429 -6348 462 -6305
rect 396 -6348 429 -6305
rect 495 -6348 528 -6305
rect 561 -6348 594 -6305
rect 594 -6348 627 -6305
rect 627 -6348 660 -6305
rect 693 -6348 726 -6305
rect 726 -6348 759 -6305
rect 759 -6348 792 -6305
rect 825 -6348 858 -6305
rect 858 -6348 891 -6305
rect 891 -6348 924 -6305
rect -33 -6419 0 -6376
rect 33 -6419 66 -6376
rect 0 -6419 33 -6376
rect 99 -6419 132 -6376
rect 165 -6419 198 -6376
rect 198 -6419 231 -6376
rect 231 -6419 264 -6376
rect 297 -6419 330 -6376
rect 264 -6419 297 -6376
rect 363 -6419 396 -6376
rect 429 -6419 462 -6376
rect 396 -6419 429 -6376
rect 495 -6419 528 -6376
rect 561 -6419 594 -6376
rect 594 -6419 627 -6376
rect 627 -6419 660 -6376
rect 693 -6419 726 -6376
rect 726 -6419 759 -6376
rect 759 -6419 792 -6376
rect 825 -6419 858 -6376
rect 792 -6419 825 -6376
rect 891 -6419 924 -6376
rect -33 -6490 0 -6447
rect 33 -6490 66 -6447
rect 0 -6490 33 -6447
rect 99 -6490 132 -6447
rect 165 -6490 198 -6447
rect 198 -6490 231 -6447
rect 231 -6490 264 -6447
rect 297 -6490 330 -6447
rect 264 -6490 297 -6447
rect 363 -6490 396 -6447
rect 429 -6490 462 -6447
rect 396 -6490 429 -6447
rect 495 -6490 528 -6447
rect 561 -6490 594 -6447
rect 594 -6490 627 -6447
rect 627 -6490 660 -6447
rect 693 -6490 726 -6447
rect 660 -6490 693 -6447
rect 759 -6490 792 -6447
rect 825 -6490 858 -6447
rect 858 -6490 891 -6447
rect 891 -6490 924 -6447
rect -33 -6561 0 -6518
rect 33 -6561 66 -6518
rect 0 -6561 33 -6518
rect 99 -6561 132 -6518
rect 165 -6561 198 -6518
rect 198 -6561 231 -6518
rect 231 -6561 264 -6518
rect 297 -6561 330 -6518
rect 264 -6561 297 -6518
rect 363 -6561 396 -6518
rect 429 -6561 462 -6518
rect 396 -6561 429 -6518
rect 495 -6561 528 -6518
rect 561 -6561 594 -6518
rect 594 -6561 627 -6518
rect 627 -6561 660 -6518
rect 693 -6561 726 -6518
rect 660 -6561 693 -6518
rect 759 -6561 792 -6518
rect 825 -6561 858 -6518
rect 792 -6561 825 -6518
rect 891 -6561 924 -6518
rect -33 -6632 0 -6589
rect 33 -6632 66 -6589
rect 0 -6632 33 -6589
rect 99 -6632 132 -6589
rect 165 -6632 198 -6589
rect 198 -6632 231 -6589
rect 231 -6632 264 -6589
rect 297 -6632 330 -6589
rect 264 -6632 297 -6589
rect 363 -6632 396 -6589
rect 429 -6632 462 -6589
rect 396 -6632 429 -6589
rect 495 -6632 528 -6589
rect 561 -6632 594 -6589
rect 528 -6632 561 -6589
rect 627 -6632 660 -6589
rect 693 -6632 726 -6589
rect 726 -6632 759 -6589
rect 759 -6632 792 -6589
rect 825 -6632 858 -6589
rect 858 -6632 891 -6589
rect 891 -6632 924 -6589
rect -33 -6703 0 -6660
rect 33 -6703 66 -6660
rect 0 -6703 33 -6660
rect 99 -6703 132 -6660
rect 165 -6703 198 -6660
rect 198 -6703 231 -6660
rect 231 -6703 264 -6660
rect 297 -6703 330 -6660
rect 264 -6703 297 -6660
rect 363 -6703 396 -6660
rect 429 -6703 462 -6660
rect 396 -6703 429 -6660
rect 495 -6703 528 -6660
rect 561 -6703 594 -6660
rect 528 -6703 561 -6660
rect 627 -6703 660 -6660
rect 693 -6703 726 -6660
rect 726 -6703 759 -6660
rect 759 -6703 792 -6660
rect 825 -6703 858 -6660
rect 792 -6703 825 -6660
rect 891 -6703 924 -6660
rect -33 -6774 0 -6731
rect 33 -6774 66 -6731
rect 0 -6774 33 -6731
rect 99 -6774 132 -6731
rect 165 -6774 198 -6731
rect 198 -6774 231 -6731
rect 231 -6774 264 -6731
rect 297 -6774 330 -6731
rect 264 -6774 297 -6731
rect 363 -6774 396 -6731
rect 429 -6774 462 -6731
rect 396 -6774 429 -6731
rect 495 -6774 528 -6731
rect 561 -6774 594 -6731
rect 528 -6774 561 -6731
rect 627 -6774 660 -6731
rect 693 -6774 726 -6731
rect 660 -6774 693 -6731
rect 759 -6774 792 -6731
rect 825 -6774 858 -6731
rect 858 -6774 891 -6731
rect 891 -6774 924 -6731
rect -33 -6845 0 -6802
rect 33 -6845 66 -6802
rect 0 -6845 33 -6802
rect 99 -6845 132 -6802
rect 165 -6845 198 -6802
rect 198 -6845 231 -6802
rect 231 -6845 264 -6802
rect 297 -6845 330 -6802
rect 264 -6845 297 -6802
rect 363 -6845 396 -6802
rect 429 -6845 462 -6802
rect 396 -6845 429 -6802
rect 495 -6845 528 -6802
rect 561 -6845 594 -6802
rect 528 -6845 561 -6802
rect 627 -6845 660 -6802
rect 693 -6845 726 -6802
rect 660 -6845 693 -6802
rect 759 -6845 792 -6802
rect 825 -6845 858 -6802
rect 792 -6845 825 -6802
rect 891 -6845 924 -6802
rect -33 -6916 0 -6873
rect 33 -6916 66 -6873
rect 0 -6916 33 -6873
rect 99 -6916 132 -6873
rect 165 -6916 198 -6873
rect 132 -6916 165 -6873
rect 231 -6916 264 -6873
rect 297 -6916 330 -6873
rect 330 -6916 363 -6873
rect 363 -6916 396 -6873
rect 429 -6916 462 -6873
rect 462 -6916 495 -6873
rect 495 -6916 528 -6873
rect 561 -6916 594 -6873
rect 594 -6916 627 -6873
rect 627 -6916 660 -6873
rect 693 -6916 726 -6873
rect 726 -6916 759 -6873
rect 759 -6916 792 -6873
rect 825 -6916 858 -6873
rect 858 -6916 891 -6873
rect 891 -6916 924 -6873
rect -33 -6987 0 -6944
rect 33 -6987 66 -6944
rect 0 -6987 33 -6944
rect 99 -6987 132 -6944
rect 165 -6987 198 -6944
rect 132 -6987 165 -6944
rect 231 -6987 264 -6944
rect 297 -6987 330 -6944
rect 330 -6987 363 -6944
rect 363 -6987 396 -6944
rect 429 -6987 462 -6944
rect 462 -6987 495 -6944
rect 495 -6987 528 -6944
rect 561 -6987 594 -6944
rect 594 -6987 627 -6944
rect 627 -6987 660 -6944
rect 693 -6987 726 -6944
rect 726 -6987 759 -6944
rect 759 -6987 792 -6944
rect 825 -6987 858 -6944
rect 792 -6987 825 -6944
rect 891 -6987 924 -6944
rect -33 -7058 0 -7015
rect 33 -7058 66 -7015
rect 0 -7058 33 -7015
rect 99 -7058 132 -7015
rect 165 -7058 198 -7015
rect 132 -7058 165 -7015
rect 231 -7058 264 -7015
rect 297 -7058 330 -7015
rect 330 -7058 363 -7015
rect 363 -7058 396 -7015
rect 429 -7058 462 -7015
rect 462 -7058 495 -7015
rect 495 -7058 528 -7015
rect 561 -7058 594 -7015
rect 594 -7058 627 -7015
rect 627 -7058 660 -7015
rect 693 -7058 726 -7015
rect 660 -7058 693 -7015
rect 759 -7058 792 -7015
rect 825 -7058 858 -7015
rect 858 -7058 891 -7015
rect 891 -7058 924 -7015
rect -33 -7129 0 -7086
rect 33 -7129 66 -7086
rect 0 -7129 33 -7086
rect 99 -7129 132 -7086
rect 165 -7129 198 -7086
rect 132 -7129 165 -7086
rect 231 -7129 264 -7086
rect 297 -7129 330 -7086
rect 330 -7129 363 -7086
rect 363 -7129 396 -7086
rect 429 -7129 462 -7086
rect 462 -7129 495 -7086
rect 495 -7129 528 -7086
rect 561 -7129 594 -7086
rect 594 -7129 627 -7086
rect 627 -7129 660 -7086
rect 693 -7129 726 -7086
rect 660 -7129 693 -7086
rect 759 -7129 792 -7086
rect 825 -7129 858 -7086
rect 792 -7129 825 -7086
rect 891 -7129 924 -7086
rect -33 -7200 0 -7157
rect 33 -7200 66 -7157
rect 0 -7200 33 -7157
rect 99 -7200 132 -7157
rect 165 -7200 198 -7157
rect 132 -7200 165 -7157
rect 231 -7200 264 -7157
rect 297 -7200 330 -7157
rect 330 -7200 363 -7157
rect 363 -7200 396 -7157
rect 429 -7200 462 -7157
rect 462 -7200 495 -7157
rect 495 -7200 528 -7157
rect 561 -7200 594 -7157
rect 528 -7200 561 -7157
rect 627 -7200 660 -7157
rect 693 -7200 726 -7157
rect 726 -7200 759 -7157
rect 759 -7200 792 -7157
rect 825 -7200 858 -7157
rect 858 -7200 891 -7157
rect 891 -7200 924 -7157
rect -33 -7271 0 -7228
rect 33 -7271 66 -7228
rect 0 -7271 33 -7228
rect 99 -7271 132 -7228
rect 165 -7271 198 -7228
rect 132 -7271 165 -7228
rect 231 -7271 264 -7228
rect 297 -7271 330 -7228
rect 330 -7271 363 -7228
rect 363 -7271 396 -7228
rect 429 -7271 462 -7228
rect 462 -7271 495 -7228
rect 495 -7271 528 -7228
rect 561 -7271 594 -7228
rect 528 -7271 561 -7228
rect 627 -7271 660 -7228
rect 693 -7271 726 -7228
rect 726 -7271 759 -7228
rect 759 -7271 792 -7228
rect 825 -7271 858 -7228
rect 792 -7271 825 -7228
rect 891 -7271 924 -7228
rect -33 -7342 0 -7299
rect 33 -7342 66 -7299
rect 0 -7342 33 -7299
rect 99 -7342 132 -7299
rect 165 -7342 198 -7299
rect 132 -7342 165 -7299
rect 231 -7342 264 -7299
rect 297 -7342 330 -7299
rect 330 -7342 363 -7299
rect 363 -7342 396 -7299
rect 429 -7342 462 -7299
rect 462 -7342 495 -7299
rect 495 -7342 528 -7299
rect 561 -7342 594 -7299
rect 528 -7342 561 -7299
rect 627 -7342 660 -7299
rect 693 -7342 726 -7299
rect 660 -7342 693 -7299
rect 759 -7342 792 -7299
rect 825 -7342 858 -7299
rect 858 -7342 891 -7299
rect 891 -7342 924 -7299
rect -33 -7413 0 -7370
rect 33 -7413 66 -7370
rect 0 -7413 33 -7370
rect 99 -7413 132 -7370
rect 165 -7413 198 -7370
rect 132 -7413 165 -7370
rect 231 -7413 264 -7370
rect 297 -7413 330 -7370
rect 330 -7413 363 -7370
rect 363 -7413 396 -7370
rect 429 -7413 462 -7370
rect 462 -7413 495 -7370
rect 495 -7413 528 -7370
rect 561 -7413 594 -7370
rect 528 -7413 561 -7370
rect 627 -7413 660 -7370
rect 693 -7413 726 -7370
rect 660 -7413 693 -7370
rect 759 -7413 792 -7370
rect 825 -7413 858 -7370
rect 792 -7413 825 -7370
rect 891 -7413 924 -7370
rect -33 -7484 0 -7441
rect 33 -7484 66 -7441
rect 0 -7484 33 -7441
rect 99 -7484 132 -7441
rect 165 -7484 198 -7441
rect 132 -7484 165 -7441
rect 231 -7484 264 -7441
rect 297 -7484 330 -7441
rect 330 -7484 363 -7441
rect 363 -7484 396 -7441
rect 429 -7484 462 -7441
rect 396 -7484 429 -7441
rect 495 -7484 528 -7441
rect 561 -7484 594 -7441
rect 594 -7484 627 -7441
rect 627 -7484 660 -7441
rect 693 -7484 726 -7441
rect 726 -7484 759 -7441
rect 759 -7484 792 -7441
rect 825 -7484 858 -7441
rect 858 -7484 891 -7441
rect 891 -7484 924 -7441
rect -33 -7555 0 -7512
rect 33 -7555 66 -7512
rect 0 -7555 33 -7512
rect 99 -7555 132 -7512
rect 165 -7555 198 -7512
rect 132 -7555 165 -7512
rect 231 -7555 264 -7512
rect 297 -7555 330 -7512
rect 330 -7555 363 -7512
rect 363 -7555 396 -7512
rect 429 -7555 462 -7512
rect 396 -7555 429 -7512
rect 495 -7555 528 -7512
rect 561 -7555 594 -7512
rect 594 -7555 627 -7512
rect 627 -7555 660 -7512
rect 693 -7555 726 -7512
rect 726 -7555 759 -7512
rect 759 -7555 792 -7512
rect 825 -7555 858 -7512
rect 792 -7555 825 -7512
rect 891 -7555 924 -7512
rect -33 -7626 0 -7583
rect 33 -7626 66 -7583
rect 0 -7626 33 -7583
rect 99 -7626 132 -7583
rect 165 -7626 198 -7583
rect 132 -7626 165 -7583
rect 231 -7626 264 -7583
rect 297 -7626 330 -7583
rect 330 -7626 363 -7583
rect 363 -7626 396 -7583
rect 429 -7626 462 -7583
rect 396 -7626 429 -7583
rect 495 -7626 528 -7583
rect 561 -7626 594 -7583
rect 594 -7626 627 -7583
rect 627 -7626 660 -7583
rect 693 -7626 726 -7583
rect 660 -7626 693 -7583
rect 759 -7626 792 -7583
rect 825 -7626 858 -7583
rect 858 -7626 891 -7583
rect 891 -7626 924 -7583
rect -33 -7697 0 -7654
rect 33 -7697 66 -7654
rect 0 -7697 33 -7654
rect 99 -7697 132 -7654
rect 165 -7697 198 -7654
rect 132 -7697 165 -7654
rect 231 -7697 264 -7654
rect 297 -7697 330 -7654
rect 330 -7697 363 -7654
rect 363 -7697 396 -7654
rect 429 -7697 462 -7654
rect 396 -7697 429 -7654
rect 495 -7697 528 -7654
rect 561 -7697 594 -7654
rect 594 -7697 627 -7654
rect 627 -7697 660 -7654
rect 693 -7697 726 -7654
rect 660 -7697 693 -7654
rect 759 -7697 792 -7654
rect 825 -7697 858 -7654
rect 792 -7697 825 -7654
rect 891 -7697 924 -7654
rect -33 -7768 0 -7725
rect 33 -7768 66 -7725
rect 0 -7768 33 -7725
rect 99 -7768 132 -7725
rect 165 -7768 198 -7725
rect 132 -7768 165 -7725
rect 231 -7768 264 -7725
rect 297 -7768 330 -7725
rect 330 -7768 363 -7725
rect 363 -7768 396 -7725
rect 429 -7768 462 -7725
rect 396 -7768 429 -7725
rect 495 -7768 528 -7725
rect 561 -7768 594 -7725
rect 528 -7768 561 -7725
rect 627 -7768 660 -7725
rect 693 -7768 726 -7725
rect 726 -7768 759 -7725
rect 759 -7768 792 -7725
rect 825 -7768 858 -7725
rect 858 -7768 891 -7725
rect 891 -7768 924 -7725
rect -33 -7839 0 -7796
rect 33 -7839 66 -7796
rect 0 -7839 33 -7796
rect 99 -7839 132 -7796
rect 165 -7839 198 -7796
rect 132 -7839 165 -7796
rect 231 -7839 264 -7796
rect 297 -7839 330 -7796
rect 330 -7839 363 -7796
rect 363 -7839 396 -7796
rect 429 -7839 462 -7796
rect 396 -7839 429 -7796
rect 495 -7839 528 -7796
rect 561 -7839 594 -7796
rect 528 -7839 561 -7796
rect 627 -7839 660 -7796
rect 693 -7839 726 -7796
rect 726 -7839 759 -7796
rect 759 -7839 792 -7796
rect 825 -7839 858 -7796
rect 792 -7839 825 -7796
rect 891 -7839 924 -7796
rect -33 -7910 0 -7867
rect 33 -7910 66 -7867
rect 0 -7910 33 -7867
rect 99 -7910 132 -7867
rect 165 -7910 198 -7867
rect 132 -7910 165 -7867
rect 231 -7910 264 -7867
rect 297 -7910 330 -7867
rect 330 -7910 363 -7867
rect 363 -7910 396 -7867
rect 429 -7910 462 -7867
rect 396 -7910 429 -7867
rect 495 -7910 528 -7867
rect 561 -7910 594 -7867
rect 528 -7910 561 -7867
rect 627 -7910 660 -7867
rect 693 -7910 726 -7867
rect 660 -7910 693 -7867
rect 759 -7910 792 -7867
rect 825 -7910 858 -7867
rect 858 -7910 891 -7867
rect 891 -7910 924 -7867
rect -33 -7981 0 -7938
rect 33 -7981 66 -7938
rect 0 -7981 33 -7938
rect 99 -7981 132 -7938
rect 165 -7981 198 -7938
rect 132 -7981 165 -7938
rect 231 -7981 264 -7938
rect 297 -7981 330 -7938
rect 330 -7981 363 -7938
rect 363 -7981 396 -7938
rect 429 -7981 462 -7938
rect 396 -7981 429 -7938
rect 495 -7981 528 -7938
rect 561 -7981 594 -7938
rect 528 -7981 561 -7938
rect 627 -7981 660 -7938
rect 693 -7981 726 -7938
rect 660 -7981 693 -7938
rect 759 -7981 792 -7938
rect 825 -7981 858 -7938
rect 792 -7981 825 -7938
rect 891 -7981 924 -7938
rect -33 -8052 0 -8009
rect 33 -8052 66 -8009
rect 0 -8052 33 -8009
rect 99 -8052 132 -8009
rect 165 -8052 198 -8009
rect 132 -8052 165 -8009
rect 231 -8052 264 -8009
rect 297 -8052 330 -8009
rect 264 -8052 297 -8009
rect 363 -8052 396 -8009
rect 429 -8052 462 -8009
rect 462 -8052 495 -8009
rect 495 -8052 528 -8009
rect 561 -8052 594 -8009
rect 594 -8052 627 -8009
rect 627 -8052 660 -8009
rect 693 -8052 726 -8009
rect 726 -8052 759 -8009
rect 759 -8052 792 -8009
rect 825 -8052 858 -8009
rect 858 -8052 891 -8009
rect 891 -8052 924 -8009
rect -33 -8123 0 -8080
rect 33 -8123 66 -8080
rect 0 -8123 33 -8080
rect 99 -8123 132 -8080
rect 165 -8123 198 -8080
rect 132 -8123 165 -8080
rect 231 -8123 264 -8080
rect 297 -8123 330 -8080
rect 264 -8123 297 -8080
rect 363 -8123 396 -8080
rect 429 -8123 462 -8080
rect 462 -8123 495 -8080
rect 495 -8123 528 -8080
rect 561 -8123 594 -8080
rect 594 -8123 627 -8080
rect 627 -8123 660 -8080
rect 693 -8123 726 -8080
rect 726 -8123 759 -8080
rect 759 -8123 792 -8080
rect 825 -8123 858 -8080
rect 792 -8123 825 -8080
rect 891 -8123 924 -8080
rect -33 -8194 0 -8151
rect 33 -8194 66 -8151
rect 0 -8194 33 -8151
rect 99 -8194 132 -8151
rect 165 -8194 198 -8151
rect 132 -8194 165 -8151
rect 231 -8194 264 -8151
rect 297 -8194 330 -8151
rect 264 -8194 297 -8151
rect 363 -8194 396 -8151
rect 429 -8194 462 -8151
rect 462 -8194 495 -8151
rect 495 -8194 528 -8151
rect 561 -8194 594 -8151
rect 594 -8194 627 -8151
rect 627 -8194 660 -8151
rect 693 -8194 726 -8151
rect 660 -8194 693 -8151
rect 759 -8194 792 -8151
rect 825 -8194 858 -8151
rect 858 -8194 891 -8151
rect 891 -8194 924 -8151
rect -33 -8265 0 -8222
rect 33 -8265 66 -8222
rect 0 -8265 33 -8222
rect 99 -8265 132 -8222
rect 165 -8265 198 -8222
rect 132 -8265 165 -8222
rect 231 -8265 264 -8222
rect 297 -8265 330 -8222
rect 264 -8265 297 -8222
rect 363 -8265 396 -8222
rect 429 -8265 462 -8222
rect 462 -8265 495 -8222
rect 495 -8265 528 -8222
rect 561 -8265 594 -8222
rect 594 -8265 627 -8222
rect 627 -8265 660 -8222
rect 693 -8265 726 -8222
rect 660 -8265 693 -8222
rect 759 -8265 792 -8222
rect 825 -8265 858 -8222
rect 792 -8265 825 -8222
rect 891 -8265 924 -8222
rect -33 -8336 0 -8293
rect 33 -8336 66 -8293
rect 0 -8336 33 -8293
rect 99 -8336 132 -8293
rect 165 -8336 198 -8293
rect 132 -8336 165 -8293
rect 231 -8336 264 -8293
rect 297 -8336 330 -8293
rect 264 -8336 297 -8293
rect 363 -8336 396 -8293
rect 429 -8336 462 -8293
rect 462 -8336 495 -8293
rect 495 -8336 528 -8293
rect 561 -8336 594 -8293
rect 528 -8336 561 -8293
rect 627 -8336 660 -8293
rect 693 -8336 726 -8293
rect 726 -8336 759 -8293
rect 759 -8336 792 -8293
rect 825 -8336 858 -8293
rect 858 -8336 891 -8293
rect 891 -8336 924 -8293
rect -33 -8407 0 -8364
rect 33 -8407 66 -8364
rect 0 -8407 33 -8364
rect 99 -8407 132 -8364
rect 165 -8407 198 -8364
rect 132 -8407 165 -8364
rect 231 -8407 264 -8364
rect 297 -8407 330 -8364
rect 264 -8407 297 -8364
rect 363 -8407 396 -8364
rect 429 -8407 462 -8364
rect 462 -8407 495 -8364
rect 495 -8407 528 -8364
rect 561 -8407 594 -8364
rect 528 -8407 561 -8364
rect 627 -8407 660 -8364
rect 693 -8407 726 -8364
rect 726 -8407 759 -8364
rect 759 -8407 792 -8364
rect 825 -8407 858 -8364
rect 792 -8407 825 -8364
rect 891 -8407 924 -8364
rect -33 -8478 0 -8435
rect 33 -8478 66 -8435
rect 0 -8478 33 -8435
rect 99 -8478 132 -8435
rect 165 -8478 198 -8435
rect 132 -8478 165 -8435
rect 231 -8478 264 -8435
rect 297 -8478 330 -8435
rect 264 -8478 297 -8435
rect 363 -8478 396 -8435
rect 429 -8478 462 -8435
rect 462 -8478 495 -8435
rect 495 -8478 528 -8435
rect 561 -8478 594 -8435
rect 528 -8478 561 -8435
rect 627 -8478 660 -8435
rect 693 -8478 726 -8435
rect 660 -8478 693 -8435
rect 759 -8478 792 -8435
rect 825 -8478 858 -8435
rect 858 -8478 891 -8435
rect 891 -8478 924 -8435
rect -33 -8549 0 -8506
rect 33 -8549 66 -8506
rect 0 -8549 33 -8506
rect 99 -8549 132 -8506
rect 165 -8549 198 -8506
rect 132 -8549 165 -8506
rect 231 -8549 264 -8506
rect 297 -8549 330 -8506
rect 264 -8549 297 -8506
rect 363 -8549 396 -8506
rect 429 -8549 462 -8506
rect 462 -8549 495 -8506
rect 495 -8549 528 -8506
rect 561 -8549 594 -8506
rect 528 -8549 561 -8506
rect 627 -8549 660 -8506
rect 693 -8549 726 -8506
rect 660 -8549 693 -8506
rect 759 -8549 792 -8506
rect 825 -8549 858 -8506
rect 792 -8549 825 -8506
rect 891 -8549 924 -8506
rect -33 -8620 0 -8577
rect 33 -8620 66 -8577
rect 0 -8620 33 -8577
rect 99 -8620 132 -8577
rect 165 -8620 198 -8577
rect 132 -8620 165 -8577
rect 231 -8620 264 -8577
rect 297 -8620 330 -8577
rect 264 -8620 297 -8577
rect 363 -8620 396 -8577
rect 429 -8620 462 -8577
rect 396 -8620 429 -8577
rect 495 -8620 528 -8577
rect 561 -8620 594 -8577
rect 594 -8620 627 -8577
rect 627 -8620 660 -8577
rect 693 -8620 726 -8577
rect 726 -8620 759 -8577
rect 759 -8620 792 -8577
rect 825 -8620 858 -8577
rect 858 -8620 891 -8577
rect 891 -8620 924 -8577
rect -33 -8691 0 -8648
rect 33 -8691 66 -8648
rect 0 -8691 33 -8648
rect 99 -8691 132 -8648
rect 165 -8691 198 -8648
rect 132 -8691 165 -8648
rect 231 -8691 264 -8648
rect 297 -8691 330 -8648
rect 264 -8691 297 -8648
rect 363 -8691 396 -8648
rect 429 -8691 462 -8648
rect 396 -8691 429 -8648
rect 495 -8691 528 -8648
rect 561 -8691 594 -8648
rect 594 -8691 627 -8648
rect 627 -8691 660 -8648
rect 693 -8691 726 -8648
rect 726 -8691 759 -8648
rect 759 -8691 792 -8648
rect 825 -8691 858 -8648
rect 792 -8691 825 -8648
rect 891 -8691 924 -8648
rect -33 -8762 0 -8719
rect 33 -8762 66 -8719
rect 0 -8762 33 -8719
rect 99 -8762 132 -8719
rect 165 -8762 198 -8719
rect 132 -8762 165 -8719
rect 231 -8762 264 -8719
rect 297 -8762 330 -8719
rect 264 -8762 297 -8719
rect 363 -8762 396 -8719
rect 429 -8762 462 -8719
rect 396 -8762 429 -8719
rect 495 -8762 528 -8719
rect 561 -8762 594 -8719
rect 594 -8762 627 -8719
rect 627 -8762 660 -8719
rect 693 -8762 726 -8719
rect 660 -8762 693 -8719
rect 759 -8762 792 -8719
rect 825 -8762 858 -8719
rect 858 -8762 891 -8719
rect 891 -8762 924 -8719
rect -33 -8833 0 -8790
rect 33 -8833 66 -8790
rect 0 -8833 33 -8790
rect 99 -8833 132 -8790
rect 165 -8833 198 -8790
rect 132 -8833 165 -8790
rect 231 -8833 264 -8790
rect 297 -8833 330 -8790
rect 264 -8833 297 -8790
rect 363 -8833 396 -8790
rect 429 -8833 462 -8790
rect 396 -8833 429 -8790
rect 495 -8833 528 -8790
rect 561 -8833 594 -8790
rect 594 -8833 627 -8790
rect 627 -8833 660 -8790
rect 693 -8833 726 -8790
rect 660 -8833 693 -8790
rect 759 -8833 792 -8790
rect 825 -8833 858 -8790
rect 792 -8833 825 -8790
rect 891 -8833 924 -8790
rect -33 -8904 0 -8861
rect 33 -8904 66 -8861
rect 0 -8904 33 -8861
rect 99 -8904 132 -8861
rect 165 -8904 198 -8861
rect 132 -8904 165 -8861
rect 231 -8904 264 -8861
rect 297 -8904 330 -8861
rect 264 -8904 297 -8861
rect 363 -8904 396 -8861
rect 429 -8904 462 -8861
rect 396 -8904 429 -8861
rect 495 -8904 528 -8861
rect 561 -8904 594 -8861
rect 528 -8904 561 -8861
rect 627 -8904 660 -8861
rect 693 -8904 726 -8861
rect 726 -8904 759 -8861
rect 759 -8904 792 -8861
rect 825 -8904 858 -8861
rect 858 -8904 891 -8861
rect 891 -8904 924 -8861
rect -33 -8975 0 -8932
rect 33 -8975 66 -8932
rect 0 -8975 33 -8932
rect 99 -8975 132 -8932
rect 165 -8975 198 -8932
rect 132 -8975 165 -8932
rect 231 -8975 264 -8932
rect 297 -8975 330 -8932
rect 264 -8975 297 -8932
rect 363 -8975 396 -8932
rect 429 -8975 462 -8932
rect 396 -8975 429 -8932
rect 495 -8975 528 -8932
rect 561 -8975 594 -8932
rect 528 -8975 561 -8932
rect 627 -8975 660 -8932
rect 693 -8975 726 -8932
rect 726 -8975 759 -8932
rect 759 -8975 792 -8932
rect 825 -8975 858 -8932
rect 792 -8975 825 -8932
rect 891 -8975 924 -8932
rect -33 -9046 0 -9003
rect 33 -9046 66 -9003
rect 0 -9046 33 -9003
rect 99 -9046 132 -9003
rect 165 -9046 198 -9003
rect 132 -9046 165 -9003
rect 231 -9046 264 -9003
rect 297 -9046 330 -9003
rect 264 -9046 297 -9003
rect 363 -9046 396 -9003
rect 429 -9046 462 -9003
rect 396 -9046 429 -9003
rect 495 -9046 528 -9003
rect 561 -9046 594 -9003
rect 528 -9046 561 -9003
rect 627 -9046 660 -9003
rect 693 -9046 726 -9003
rect 660 -9046 693 -9003
rect 759 -9046 792 -9003
rect 825 -9046 858 -9003
rect 858 -9046 891 -9003
rect 891 -9046 924 -9003
rect -33 -9117 0 -9074
rect 33 -9117 66 -9074
rect 0 -9117 33 -9074
rect 99 -9117 132 -9074
rect 165 -9117 198 -9074
rect 132 -9117 165 -9074
rect 231 -9117 264 -9074
rect 297 -9117 330 -9074
rect 264 -9117 297 -9074
rect 363 -9117 396 -9074
rect 429 -9117 462 -9074
rect 396 -9117 429 -9074
rect 495 -9117 528 -9074
rect 561 -9117 594 -9074
rect 528 -9117 561 -9074
rect 627 -9117 660 -9074
rect 693 -9117 726 -9074
rect 660 -9117 693 -9074
rect 759 -9117 792 -9074
rect 825 -9117 858 -9074
rect 792 -9117 825 -9074
rect 891 -9117 924 -9074
rect 56 82 89 125
rect 0 82 56 125
rect 188 82 221 125
rect 132 82 188 125
rect 320 82 353 125
rect 264 82 320 125
rect 452 82 485 125
rect 396 82 452 125
rect 584 82 617 125
rect 528 82 584 125
rect 716 82 749 125
rect 660 82 716 125
rect 848 82 881 125
rect 792 82 848 125
rect 1065 82 1098 125
rect 1098 82 1154 125
rect 1197 82 1230 125
rect 1230 82 1286 125
rect 1329 82 1362 125
rect 1362 82 1418 125
rect 1461 82 1494 125
rect 1494 82 1550 125
rect 1593 82 1626 125
rect 1626 82 1682 125
rect 1725 82 1758 125
rect 1758 82 1814 125
rect 1857 82 1890 125
rect 1890 82 1946 125
<< ndiff >>
rect 1022 -100 1055 -57
rect 1055 -100 1088 -57
rect 1088 -100 1121 -57
rect 1154 -100 1187 -57
rect 1187 -100 1220 -57
rect 1220 -100 1253 -57
rect 1286 -100 1319 -57
rect 1319 -100 1352 -57
rect 1352 -100 1385 -57
rect 1418 -100 1451 -57
rect 1451 -100 1484 -57
rect 1484 -100 1517 -57
rect 1550 -100 1583 -57
rect 1583 -100 1616 -57
rect 1616 -100 1649 -57
rect 1682 -100 1715 -57
rect 1715 -100 1748 -57
rect 1748 -100 1781 -57
rect 1814 -100 1847 -57
rect 1847 -100 1880 -57
rect 1880 -100 1913 -57
rect 1121 -171 1154 -128
rect 1154 -171 1187 -128
rect 1088 -171 1121 -128
rect 1154 -171 1187 -128
rect 1187 -171 1220 -128
rect 1220 -171 1253 -128
rect 1286 -171 1319 -128
rect 1319 -171 1352 -128
rect 1352 -171 1385 -128
rect 1418 -171 1451 -128
rect 1451 -171 1484 -128
rect 1484 -171 1517 -128
rect 1550 -171 1583 -128
rect 1583 -171 1616 -128
rect 1616 -171 1649 -128
rect 1682 -171 1715 -128
rect 1715 -171 1748 -128
rect 1748 -171 1781 -128
rect 1814 -171 1847 -128
rect 1847 -171 1880 -128
rect 1880 -171 1913 -128
rect 1022 -242 1055 -199
rect 1055 -242 1088 -199
rect 1088 -242 1121 -199
rect 1253 -242 1286 -199
rect 1286 -242 1319 -199
rect 1220 -242 1253 -199
rect 1286 -242 1319 -199
rect 1319 -242 1352 -199
rect 1352 -242 1385 -199
rect 1418 -242 1451 -199
rect 1451 -242 1484 -199
rect 1484 -242 1517 -199
rect 1550 -242 1583 -199
rect 1583 -242 1616 -199
rect 1616 -242 1649 -199
rect 1682 -242 1715 -199
rect 1715 -242 1748 -199
rect 1748 -242 1781 -199
rect 1814 -242 1847 -199
rect 1847 -242 1880 -199
rect 1880 -242 1913 -199
rect 1121 -313 1154 -270
rect 1154 -313 1187 -270
rect 1088 -313 1121 -270
rect 1253 -313 1286 -270
rect 1286 -313 1319 -270
rect 1220 -313 1253 -270
rect 1286 -313 1319 -270
rect 1319 -313 1352 -270
rect 1352 -313 1385 -270
rect 1418 -313 1451 -270
rect 1451 -313 1484 -270
rect 1484 -313 1517 -270
rect 1550 -313 1583 -270
rect 1583 -313 1616 -270
rect 1616 -313 1649 -270
rect 1682 -313 1715 -270
rect 1715 -313 1748 -270
rect 1748 -313 1781 -270
rect 1814 -313 1847 -270
rect 1847 -313 1880 -270
rect 1880 -313 1913 -270
rect 1022 -384 1055 -341
rect 1055 -384 1088 -341
rect 1088 -384 1121 -341
rect 1154 -384 1187 -341
rect 1187 -384 1220 -341
rect 1220 -384 1253 -341
rect 1385 -384 1418 -341
rect 1418 -384 1451 -341
rect 1352 -384 1385 -341
rect 1418 -384 1451 -341
rect 1451 -384 1484 -341
rect 1484 -384 1517 -341
rect 1550 -384 1583 -341
rect 1583 -384 1616 -341
rect 1616 -384 1649 -341
rect 1682 -384 1715 -341
rect 1715 -384 1748 -341
rect 1748 -384 1781 -341
rect 1814 -384 1847 -341
rect 1847 -384 1880 -341
rect 1880 -384 1913 -341
rect 1121 -455 1154 -412
rect 1154 -455 1187 -412
rect 1088 -455 1121 -412
rect 1154 -455 1187 -412
rect 1187 -455 1220 -412
rect 1220 -455 1253 -412
rect 1385 -455 1418 -412
rect 1418 -455 1451 -412
rect 1352 -455 1385 -412
rect 1418 -455 1451 -412
rect 1451 -455 1484 -412
rect 1484 -455 1517 -412
rect 1550 -455 1583 -412
rect 1583 -455 1616 -412
rect 1616 -455 1649 -412
rect 1682 -455 1715 -412
rect 1715 -455 1748 -412
rect 1748 -455 1781 -412
rect 1814 -455 1847 -412
rect 1847 -455 1880 -412
rect 1880 -455 1913 -412
rect 1022 -526 1055 -483
rect 1055 -526 1088 -483
rect 1088 -526 1121 -483
rect 1253 -526 1286 -483
rect 1286 -526 1319 -483
rect 1220 -526 1253 -483
rect 1385 -526 1418 -483
rect 1418 -526 1451 -483
rect 1352 -526 1385 -483
rect 1418 -526 1451 -483
rect 1451 -526 1484 -483
rect 1484 -526 1517 -483
rect 1550 -526 1583 -483
rect 1583 -526 1616 -483
rect 1616 -526 1649 -483
rect 1682 -526 1715 -483
rect 1715 -526 1748 -483
rect 1748 -526 1781 -483
rect 1814 -526 1847 -483
rect 1847 -526 1880 -483
rect 1880 -526 1913 -483
rect 1121 -597 1154 -554
rect 1154 -597 1187 -554
rect 1088 -597 1121 -554
rect 1253 -597 1286 -554
rect 1286 -597 1319 -554
rect 1220 -597 1253 -554
rect 1385 -597 1418 -554
rect 1418 -597 1451 -554
rect 1352 -597 1385 -554
rect 1418 -597 1451 -554
rect 1451 -597 1484 -554
rect 1484 -597 1517 -554
rect 1550 -597 1583 -554
rect 1583 -597 1616 -554
rect 1616 -597 1649 -554
rect 1682 -597 1715 -554
rect 1715 -597 1748 -554
rect 1748 -597 1781 -554
rect 1814 -597 1847 -554
rect 1847 -597 1880 -554
rect 1880 -597 1913 -554
rect 1022 -668 1055 -625
rect 1055 -668 1088 -625
rect 1088 -668 1121 -625
rect 1154 -668 1187 -625
rect 1187 -668 1220 -625
rect 1220 -668 1253 -625
rect 1286 -668 1319 -625
rect 1319 -668 1352 -625
rect 1352 -668 1385 -625
rect 1517 -668 1550 -625
rect 1550 -668 1583 -625
rect 1484 -668 1517 -625
rect 1550 -668 1583 -625
rect 1583 -668 1616 -625
rect 1616 -668 1649 -625
rect 1682 -668 1715 -625
rect 1715 -668 1748 -625
rect 1748 -668 1781 -625
rect 1814 -668 1847 -625
rect 1847 -668 1880 -625
rect 1880 -668 1913 -625
rect 1121 -739 1154 -696
rect 1154 -739 1187 -696
rect 1088 -739 1121 -696
rect 1154 -739 1187 -696
rect 1187 -739 1220 -696
rect 1220 -739 1253 -696
rect 1286 -739 1319 -696
rect 1319 -739 1352 -696
rect 1352 -739 1385 -696
rect 1517 -739 1550 -696
rect 1550 -739 1583 -696
rect 1484 -739 1517 -696
rect 1550 -739 1583 -696
rect 1583 -739 1616 -696
rect 1616 -739 1649 -696
rect 1682 -739 1715 -696
rect 1715 -739 1748 -696
rect 1748 -739 1781 -696
rect 1814 -739 1847 -696
rect 1847 -739 1880 -696
rect 1880 -739 1913 -696
rect 1022 -810 1055 -767
rect 1055 -810 1088 -767
rect 1088 -810 1121 -767
rect 1253 -810 1286 -767
rect 1286 -810 1319 -767
rect 1220 -810 1253 -767
rect 1286 -810 1319 -767
rect 1319 -810 1352 -767
rect 1352 -810 1385 -767
rect 1517 -810 1550 -767
rect 1550 -810 1583 -767
rect 1484 -810 1517 -767
rect 1550 -810 1583 -767
rect 1583 -810 1616 -767
rect 1616 -810 1649 -767
rect 1682 -810 1715 -767
rect 1715 -810 1748 -767
rect 1748 -810 1781 -767
rect 1814 -810 1847 -767
rect 1847 -810 1880 -767
rect 1880 -810 1913 -767
rect 1121 -881 1154 -838
rect 1154 -881 1187 -838
rect 1088 -881 1121 -838
rect 1253 -881 1286 -838
rect 1286 -881 1319 -838
rect 1220 -881 1253 -838
rect 1286 -881 1319 -838
rect 1319 -881 1352 -838
rect 1352 -881 1385 -838
rect 1517 -881 1550 -838
rect 1550 -881 1583 -838
rect 1484 -881 1517 -838
rect 1550 -881 1583 -838
rect 1583 -881 1616 -838
rect 1616 -881 1649 -838
rect 1682 -881 1715 -838
rect 1715 -881 1748 -838
rect 1748 -881 1781 -838
rect 1814 -881 1847 -838
rect 1847 -881 1880 -838
rect 1880 -881 1913 -838
rect 1022 -952 1055 -909
rect 1055 -952 1088 -909
rect 1088 -952 1121 -909
rect 1154 -952 1187 -909
rect 1187 -952 1220 -909
rect 1220 -952 1253 -909
rect 1385 -952 1418 -909
rect 1418 -952 1451 -909
rect 1352 -952 1385 -909
rect 1517 -952 1550 -909
rect 1550 -952 1583 -909
rect 1484 -952 1517 -909
rect 1550 -952 1583 -909
rect 1583 -952 1616 -909
rect 1616 -952 1649 -909
rect 1682 -952 1715 -909
rect 1715 -952 1748 -909
rect 1748 -952 1781 -909
rect 1814 -952 1847 -909
rect 1847 -952 1880 -909
rect 1880 -952 1913 -909
rect 1121 -1023 1154 -980
rect 1154 -1023 1187 -980
rect 1088 -1023 1121 -980
rect 1154 -1023 1187 -980
rect 1187 -1023 1220 -980
rect 1220 -1023 1253 -980
rect 1385 -1023 1418 -980
rect 1418 -1023 1451 -980
rect 1352 -1023 1385 -980
rect 1517 -1023 1550 -980
rect 1550 -1023 1583 -980
rect 1484 -1023 1517 -980
rect 1550 -1023 1583 -980
rect 1583 -1023 1616 -980
rect 1616 -1023 1649 -980
rect 1682 -1023 1715 -980
rect 1715 -1023 1748 -980
rect 1748 -1023 1781 -980
rect 1814 -1023 1847 -980
rect 1847 -1023 1880 -980
rect 1880 -1023 1913 -980
rect 1022 -1094 1055 -1051
rect 1055 -1094 1088 -1051
rect 1088 -1094 1121 -1051
rect 1253 -1094 1286 -1051
rect 1286 -1094 1319 -1051
rect 1220 -1094 1253 -1051
rect 1385 -1094 1418 -1051
rect 1418 -1094 1451 -1051
rect 1352 -1094 1385 -1051
rect 1517 -1094 1550 -1051
rect 1550 -1094 1583 -1051
rect 1484 -1094 1517 -1051
rect 1550 -1094 1583 -1051
rect 1583 -1094 1616 -1051
rect 1616 -1094 1649 -1051
rect 1682 -1094 1715 -1051
rect 1715 -1094 1748 -1051
rect 1748 -1094 1781 -1051
rect 1814 -1094 1847 -1051
rect 1847 -1094 1880 -1051
rect 1880 -1094 1913 -1051
rect 1121 -1165 1154 -1122
rect 1154 -1165 1187 -1122
rect 1088 -1165 1121 -1122
rect 1253 -1165 1286 -1122
rect 1286 -1165 1319 -1122
rect 1220 -1165 1253 -1122
rect 1385 -1165 1418 -1122
rect 1418 -1165 1451 -1122
rect 1352 -1165 1385 -1122
rect 1517 -1165 1550 -1122
rect 1550 -1165 1583 -1122
rect 1484 -1165 1517 -1122
rect 1550 -1165 1583 -1122
rect 1583 -1165 1616 -1122
rect 1616 -1165 1649 -1122
rect 1682 -1165 1715 -1122
rect 1715 -1165 1748 -1122
rect 1748 -1165 1781 -1122
rect 1814 -1165 1847 -1122
rect 1847 -1165 1880 -1122
rect 1880 -1165 1913 -1122
rect 1022 -1236 1055 -1193
rect 1055 -1236 1088 -1193
rect 1088 -1236 1121 -1193
rect 1154 -1236 1187 -1193
rect 1187 -1236 1220 -1193
rect 1220 -1236 1253 -1193
rect 1286 -1236 1319 -1193
rect 1319 -1236 1352 -1193
rect 1352 -1236 1385 -1193
rect 1418 -1236 1451 -1193
rect 1451 -1236 1484 -1193
rect 1484 -1236 1517 -1193
rect 1649 -1236 1682 -1193
rect 1682 -1236 1715 -1193
rect 1616 -1236 1649 -1193
rect 1682 -1236 1715 -1193
rect 1715 -1236 1748 -1193
rect 1748 -1236 1781 -1193
rect 1814 -1236 1847 -1193
rect 1847 -1236 1880 -1193
rect 1880 -1236 1913 -1193
rect 1121 -1307 1154 -1264
rect 1154 -1307 1187 -1264
rect 1088 -1307 1121 -1264
rect 1154 -1307 1187 -1264
rect 1187 -1307 1220 -1264
rect 1220 -1307 1253 -1264
rect 1286 -1307 1319 -1264
rect 1319 -1307 1352 -1264
rect 1352 -1307 1385 -1264
rect 1418 -1307 1451 -1264
rect 1451 -1307 1484 -1264
rect 1484 -1307 1517 -1264
rect 1649 -1307 1682 -1264
rect 1682 -1307 1715 -1264
rect 1616 -1307 1649 -1264
rect 1682 -1307 1715 -1264
rect 1715 -1307 1748 -1264
rect 1748 -1307 1781 -1264
rect 1814 -1307 1847 -1264
rect 1847 -1307 1880 -1264
rect 1880 -1307 1913 -1264
rect 1022 -1378 1055 -1335
rect 1055 -1378 1088 -1335
rect 1088 -1378 1121 -1335
rect 1253 -1378 1286 -1335
rect 1286 -1378 1319 -1335
rect 1220 -1378 1253 -1335
rect 1286 -1378 1319 -1335
rect 1319 -1378 1352 -1335
rect 1352 -1378 1385 -1335
rect 1418 -1378 1451 -1335
rect 1451 -1378 1484 -1335
rect 1484 -1378 1517 -1335
rect 1649 -1378 1682 -1335
rect 1682 -1378 1715 -1335
rect 1616 -1378 1649 -1335
rect 1682 -1378 1715 -1335
rect 1715 -1378 1748 -1335
rect 1748 -1378 1781 -1335
rect 1814 -1378 1847 -1335
rect 1847 -1378 1880 -1335
rect 1880 -1378 1913 -1335
rect 1121 -1449 1154 -1406
rect 1154 -1449 1187 -1406
rect 1088 -1449 1121 -1406
rect 1253 -1449 1286 -1406
rect 1286 -1449 1319 -1406
rect 1220 -1449 1253 -1406
rect 1286 -1449 1319 -1406
rect 1319 -1449 1352 -1406
rect 1352 -1449 1385 -1406
rect 1418 -1449 1451 -1406
rect 1451 -1449 1484 -1406
rect 1484 -1449 1517 -1406
rect 1649 -1449 1682 -1406
rect 1682 -1449 1715 -1406
rect 1616 -1449 1649 -1406
rect 1682 -1449 1715 -1406
rect 1715 -1449 1748 -1406
rect 1748 -1449 1781 -1406
rect 1814 -1449 1847 -1406
rect 1847 -1449 1880 -1406
rect 1880 -1449 1913 -1406
rect 1022 -1520 1055 -1477
rect 1055 -1520 1088 -1477
rect 1088 -1520 1121 -1477
rect 1154 -1520 1187 -1477
rect 1187 -1520 1220 -1477
rect 1220 -1520 1253 -1477
rect 1385 -1520 1418 -1477
rect 1418 -1520 1451 -1477
rect 1352 -1520 1385 -1477
rect 1418 -1520 1451 -1477
rect 1451 -1520 1484 -1477
rect 1484 -1520 1517 -1477
rect 1649 -1520 1682 -1477
rect 1682 -1520 1715 -1477
rect 1616 -1520 1649 -1477
rect 1682 -1520 1715 -1477
rect 1715 -1520 1748 -1477
rect 1748 -1520 1781 -1477
rect 1814 -1520 1847 -1477
rect 1847 -1520 1880 -1477
rect 1880 -1520 1913 -1477
rect 1121 -1591 1154 -1548
rect 1154 -1591 1187 -1548
rect 1088 -1591 1121 -1548
rect 1154 -1591 1187 -1548
rect 1187 -1591 1220 -1548
rect 1220 -1591 1253 -1548
rect 1385 -1591 1418 -1548
rect 1418 -1591 1451 -1548
rect 1352 -1591 1385 -1548
rect 1418 -1591 1451 -1548
rect 1451 -1591 1484 -1548
rect 1484 -1591 1517 -1548
rect 1649 -1591 1682 -1548
rect 1682 -1591 1715 -1548
rect 1616 -1591 1649 -1548
rect 1682 -1591 1715 -1548
rect 1715 -1591 1748 -1548
rect 1748 -1591 1781 -1548
rect 1814 -1591 1847 -1548
rect 1847 -1591 1880 -1548
rect 1880 -1591 1913 -1548
rect 1022 -1662 1055 -1619
rect 1055 -1662 1088 -1619
rect 1088 -1662 1121 -1619
rect 1253 -1662 1286 -1619
rect 1286 -1662 1319 -1619
rect 1220 -1662 1253 -1619
rect 1385 -1662 1418 -1619
rect 1418 -1662 1451 -1619
rect 1352 -1662 1385 -1619
rect 1418 -1662 1451 -1619
rect 1451 -1662 1484 -1619
rect 1484 -1662 1517 -1619
rect 1649 -1662 1682 -1619
rect 1682 -1662 1715 -1619
rect 1616 -1662 1649 -1619
rect 1682 -1662 1715 -1619
rect 1715 -1662 1748 -1619
rect 1748 -1662 1781 -1619
rect 1814 -1662 1847 -1619
rect 1847 -1662 1880 -1619
rect 1880 -1662 1913 -1619
rect 1121 -1733 1154 -1690
rect 1154 -1733 1187 -1690
rect 1088 -1733 1121 -1690
rect 1253 -1733 1286 -1690
rect 1286 -1733 1319 -1690
rect 1220 -1733 1253 -1690
rect 1385 -1733 1418 -1690
rect 1418 -1733 1451 -1690
rect 1352 -1733 1385 -1690
rect 1418 -1733 1451 -1690
rect 1451 -1733 1484 -1690
rect 1484 -1733 1517 -1690
rect 1649 -1733 1682 -1690
rect 1682 -1733 1715 -1690
rect 1616 -1733 1649 -1690
rect 1682 -1733 1715 -1690
rect 1715 -1733 1748 -1690
rect 1748 -1733 1781 -1690
rect 1814 -1733 1847 -1690
rect 1847 -1733 1880 -1690
rect 1880 -1733 1913 -1690
rect 1022 -1804 1055 -1761
rect 1055 -1804 1088 -1761
rect 1088 -1804 1121 -1761
rect 1154 -1804 1187 -1761
rect 1187 -1804 1220 -1761
rect 1220 -1804 1253 -1761
rect 1286 -1804 1319 -1761
rect 1319 -1804 1352 -1761
rect 1352 -1804 1385 -1761
rect 1517 -1804 1550 -1761
rect 1550 -1804 1583 -1761
rect 1484 -1804 1517 -1761
rect 1649 -1804 1682 -1761
rect 1682 -1804 1715 -1761
rect 1616 -1804 1649 -1761
rect 1682 -1804 1715 -1761
rect 1715 -1804 1748 -1761
rect 1748 -1804 1781 -1761
rect 1814 -1804 1847 -1761
rect 1847 -1804 1880 -1761
rect 1880 -1804 1913 -1761
rect 1121 -1875 1154 -1832
rect 1154 -1875 1187 -1832
rect 1088 -1875 1121 -1832
rect 1154 -1875 1187 -1832
rect 1187 -1875 1220 -1832
rect 1220 -1875 1253 -1832
rect 1286 -1875 1319 -1832
rect 1319 -1875 1352 -1832
rect 1352 -1875 1385 -1832
rect 1517 -1875 1550 -1832
rect 1550 -1875 1583 -1832
rect 1484 -1875 1517 -1832
rect 1649 -1875 1682 -1832
rect 1682 -1875 1715 -1832
rect 1616 -1875 1649 -1832
rect 1682 -1875 1715 -1832
rect 1715 -1875 1748 -1832
rect 1748 -1875 1781 -1832
rect 1814 -1875 1847 -1832
rect 1847 -1875 1880 -1832
rect 1880 -1875 1913 -1832
rect 1022 -1946 1055 -1903
rect 1055 -1946 1088 -1903
rect 1088 -1946 1121 -1903
rect 1253 -1946 1286 -1903
rect 1286 -1946 1319 -1903
rect 1220 -1946 1253 -1903
rect 1286 -1946 1319 -1903
rect 1319 -1946 1352 -1903
rect 1352 -1946 1385 -1903
rect 1517 -1946 1550 -1903
rect 1550 -1946 1583 -1903
rect 1484 -1946 1517 -1903
rect 1649 -1946 1682 -1903
rect 1682 -1946 1715 -1903
rect 1616 -1946 1649 -1903
rect 1682 -1946 1715 -1903
rect 1715 -1946 1748 -1903
rect 1748 -1946 1781 -1903
rect 1814 -1946 1847 -1903
rect 1847 -1946 1880 -1903
rect 1880 -1946 1913 -1903
rect 1121 -2017 1154 -1974
rect 1154 -2017 1187 -1974
rect 1088 -2017 1121 -1974
rect 1253 -2017 1286 -1974
rect 1286 -2017 1319 -1974
rect 1220 -2017 1253 -1974
rect 1286 -2017 1319 -1974
rect 1319 -2017 1352 -1974
rect 1352 -2017 1385 -1974
rect 1517 -2017 1550 -1974
rect 1550 -2017 1583 -1974
rect 1484 -2017 1517 -1974
rect 1649 -2017 1682 -1974
rect 1682 -2017 1715 -1974
rect 1616 -2017 1649 -1974
rect 1682 -2017 1715 -1974
rect 1715 -2017 1748 -1974
rect 1748 -2017 1781 -1974
rect 1814 -2017 1847 -1974
rect 1847 -2017 1880 -1974
rect 1880 -2017 1913 -1974
rect 1022 -2088 1055 -2045
rect 1055 -2088 1088 -2045
rect 1088 -2088 1121 -2045
rect 1154 -2088 1187 -2045
rect 1187 -2088 1220 -2045
rect 1220 -2088 1253 -2045
rect 1385 -2088 1418 -2045
rect 1418 -2088 1451 -2045
rect 1352 -2088 1385 -2045
rect 1517 -2088 1550 -2045
rect 1550 -2088 1583 -2045
rect 1484 -2088 1517 -2045
rect 1649 -2088 1682 -2045
rect 1682 -2088 1715 -2045
rect 1616 -2088 1649 -2045
rect 1682 -2088 1715 -2045
rect 1715 -2088 1748 -2045
rect 1748 -2088 1781 -2045
rect 1814 -2088 1847 -2045
rect 1847 -2088 1880 -2045
rect 1880 -2088 1913 -2045
rect 1121 -2159 1154 -2116
rect 1154 -2159 1187 -2116
rect 1088 -2159 1121 -2116
rect 1154 -2159 1187 -2116
rect 1187 -2159 1220 -2116
rect 1220 -2159 1253 -2116
rect 1385 -2159 1418 -2116
rect 1418 -2159 1451 -2116
rect 1352 -2159 1385 -2116
rect 1517 -2159 1550 -2116
rect 1550 -2159 1583 -2116
rect 1484 -2159 1517 -2116
rect 1649 -2159 1682 -2116
rect 1682 -2159 1715 -2116
rect 1616 -2159 1649 -2116
rect 1682 -2159 1715 -2116
rect 1715 -2159 1748 -2116
rect 1748 -2159 1781 -2116
rect 1814 -2159 1847 -2116
rect 1847 -2159 1880 -2116
rect 1880 -2159 1913 -2116
rect 1022 -2230 1055 -2187
rect 1055 -2230 1088 -2187
rect 1088 -2230 1121 -2187
rect 1253 -2230 1286 -2187
rect 1286 -2230 1319 -2187
rect 1220 -2230 1253 -2187
rect 1385 -2230 1418 -2187
rect 1418 -2230 1451 -2187
rect 1352 -2230 1385 -2187
rect 1517 -2230 1550 -2187
rect 1550 -2230 1583 -2187
rect 1484 -2230 1517 -2187
rect 1649 -2230 1682 -2187
rect 1682 -2230 1715 -2187
rect 1616 -2230 1649 -2187
rect 1682 -2230 1715 -2187
rect 1715 -2230 1748 -2187
rect 1748 -2230 1781 -2187
rect 1814 -2230 1847 -2187
rect 1847 -2230 1880 -2187
rect 1880 -2230 1913 -2187
rect 1121 -2301 1154 -2258
rect 1154 -2301 1187 -2258
rect 1088 -2301 1121 -2258
rect 1253 -2301 1286 -2258
rect 1286 -2301 1319 -2258
rect 1220 -2301 1253 -2258
rect 1385 -2301 1418 -2258
rect 1418 -2301 1451 -2258
rect 1352 -2301 1385 -2258
rect 1517 -2301 1550 -2258
rect 1550 -2301 1583 -2258
rect 1484 -2301 1517 -2258
rect 1649 -2301 1682 -2258
rect 1682 -2301 1715 -2258
rect 1616 -2301 1649 -2258
rect 1682 -2301 1715 -2258
rect 1715 -2301 1748 -2258
rect 1748 -2301 1781 -2258
rect 1814 -2301 1847 -2258
rect 1847 -2301 1880 -2258
rect 1880 -2301 1913 -2258
rect 1022 -2372 1055 -2329
rect 1055 -2372 1088 -2329
rect 1088 -2372 1121 -2329
rect 1154 -2372 1187 -2329
rect 1187 -2372 1220 -2329
rect 1220 -2372 1253 -2329
rect 1286 -2372 1319 -2329
rect 1319 -2372 1352 -2329
rect 1352 -2372 1385 -2329
rect 1418 -2372 1451 -2329
rect 1451 -2372 1484 -2329
rect 1484 -2372 1517 -2329
rect 1550 -2372 1583 -2329
rect 1583 -2372 1616 -2329
rect 1616 -2372 1649 -2329
rect 1781 -2372 1814 -2329
rect 1814 -2372 1847 -2329
rect 1748 -2372 1781 -2329
rect 1814 -2372 1847 -2329
rect 1847 -2372 1880 -2329
rect 1880 -2372 1913 -2329
rect 1121 -2443 1154 -2400
rect 1154 -2443 1187 -2400
rect 1088 -2443 1121 -2400
rect 1154 -2443 1187 -2400
rect 1187 -2443 1220 -2400
rect 1220 -2443 1253 -2400
rect 1286 -2443 1319 -2400
rect 1319 -2443 1352 -2400
rect 1352 -2443 1385 -2400
rect 1418 -2443 1451 -2400
rect 1451 -2443 1484 -2400
rect 1484 -2443 1517 -2400
rect 1550 -2443 1583 -2400
rect 1583 -2443 1616 -2400
rect 1616 -2443 1649 -2400
rect 1781 -2443 1814 -2400
rect 1814 -2443 1847 -2400
rect 1748 -2443 1781 -2400
rect 1814 -2443 1847 -2400
rect 1847 -2443 1880 -2400
rect 1880 -2443 1913 -2400
rect 1022 -2514 1055 -2471
rect 1055 -2514 1088 -2471
rect 1088 -2514 1121 -2471
rect 1253 -2514 1286 -2471
rect 1286 -2514 1319 -2471
rect 1220 -2514 1253 -2471
rect 1286 -2514 1319 -2471
rect 1319 -2514 1352 -2471
rect 1352 -2514 1385 -2471
rect 1418 -2514 1451 -2471
rect 1451 -2514 1484 -2471
rect 1484 -2514 1517 -2471
rect 1550 -2514 1583 -2471
rect 1583 -2514 1616 -2471
rect 1616 -2514 1649 -2471
rect 1781 -2514 1814 -2471
rect 1814 -2514 1847 -2471
rect 1748 -2514 1781 -2471
rect 1814 -2514 1847 -2471
rect 1847 -2514 1880 -2471
rect 1880 -2514 1913 -2471
rect 1121 -2585 1154 -2542
rect 1154 -2585 1187 -2542
rect 1088 -2585 1121 -2542
rect 1253 -2585 1286 -2542
rect 1286 -2585 1319 -2542
rect 1220 -2585 1253 -2542
rect 1286 -2585 1319 -2542
rect 1319 -2585 1352 -2542
rect 1352 -2585 1385 -2542
rect 1418 -2585 1451 -2542
rect 1451 -2585 1484 -2542
rect 1484 -2585 1517 -2542
rect 1550 -2585 1583 -2542
rect 1583 -2585 1616 -2542
rect 1616 -2585 1649 -2542
rect 1781 -2585 1814 -2542
rect 1814 -2585 1847 -2542
rect 1748 -2585 1781 -2542
rect 1814 -2585 1847 -2542
rect 1847 -2585 1880 -2542
rect 1880 -2585 1913 -2542
rect 1022 -2656 1055 -2613
rect 1055 -2656 1088 -2613
rect 1088 -2656 1121 -2613
rect 1154 -2656 1187 -2613
rect 1187 -2656 1220 -2613
rect 1220 -2656 1253 -2613
rect 1385 -2656 1418 -2613
rect 1418 -2656 1451 -2613
rect 1352 -2656 1385 -2613
rect 1418 -2656 1451 -2613
rect 1451 -2656 1484 -2613
rect 1484 -2656 1517 -2613
rect 1550 -2656 1583 -2613
rect 1583 -2656 1616 -2613
rect 1616 -2656 1649 -2613
rect 1781 -2656 1814 -2613
rect 1814 -2656 1847 -2613
rect 1748 -2656 1781 -2613
rect 1814 -2656 1847 -2613
rect 1847 -2656 1880 -2613
rect 1880 -2656 1913 -2613
rect 1121 -2727 1154 -2684
rect 1154 -2727 1187 -2684
rect 1088 -2727 1121 -2684
rect 1154 -2727 1187 -2684
rect 1187 -2727 1220 -2684
rect 1220 -2727 1253 -2684
rect 1385 -2727 1418 -2684
rect 1418 -2727 1451 -2684
rect 1352 -2727 1385 -2684
rect 1418 -2727 1451 -2684
rect 1451 -2727 1484 -2684
rect 1484 -2727 1517 -2684
rect 1550 -2727 1583 -2684
rect 1583 -2727 1616 -2684
rect 1616 -2727 1649 -2684
rect 1781 -2727 1814 -2684
rect 1814 -2727 1847 -2684
rect 1748 -2727 1781 -2684
rect 1814 -2727 1847 -2684
rect 1847 -2727 1880 -2684
rect 1880 -2727 1913 -2684
rect 1022 -2798 1055 -2755
rect 1055 -2798 1088 -2755
rect 1088 -2798 1121 -2755
rect 1253 -2798 1286 -2755
rect 1286 -2798 1319 -2755
rect 1220 -2798 1253 -2755
rect 1385 -2798 1418 -2755
rect 1418 -2798 1451 -2755
rect 1352 -2798 1385 -2755
rect 1418 -2798 1451 -2755
rect 1451 -2798 1484 -2755
rect 1484 -2798 1517 -2755
rect 1550 -2798 1583 -2755
rect 1583 -2798 1616 -2755
rect 1616 -2798 1649 -2755
rect 1781 -2798 1814 -2755
rect 1814 -2798 1847 -2755
rect 1748 -2798 1781 -2755
rect 1814 -2798 1847 -2755
rect 1847 -2798 1880 -2755
rect 1880 -2798 1913 -2755
rect 1121 -2869 1154 -2826
rect 1154 -2869 1187 -2826
rect 1088 -2869 1121 -2826
rect 1253 -2869 1286 -2826
rect 1286 -2869 1319 -2826
rect 1220 -2869 1253 -2826
rect 1385 -2869 1418 -2826
rect 1418 -2869 1451 -2826
rect 1352 -2869 1385 -2826
rect 1418 -2869 1451 -2826
rect 1451 -2869 1484 -2826
rect 1484 -2869 1517 -2826
rect 1550 -2869 1583 -2826
rect 1583 -2869 1616 -2826
rect 1616 -2869 1649 -2826
rect 1781 -2869 1814 -2826
rect 1814 -2869 1847 -2826
rect 1748 -2869 1781 -2826
rect 1814 -2869 1847 -2826
rect 1847 -2869 1880 -2826
rect 1880 -2869 1913 -2826
rect 1022 -2940 1055 -2897
rect 1055 -2940 1088 -2897
rect 1088 -2940 1121 -2897
rect 1154 -2940 1187 -2897
rect 1187 -2940 1220 -2897
rect 1220 -2940 1253 -2897
rect 1286 -2940 1319 -2897
rect 1319 -2940 1352 -2897
rect 1352 -2940 1385 -2897
rect 1517 -2940 1550 -2897
rect 1550 -2940 1583 -2897
rect 1484 -2940 1517 -2897
rect 1550 -2940 1583 -2897
rect 1583 -2940 1616 -2897
rect 1616 -2940 1649 -2897
rect 1781 -2940 1814 -2897
rect 1814 -2940 1847 -2897
rect 1748 -2940 1781 -2897
rect 1814 -2940 1847 -2897
rect 1847 -2940 1880 -2897
rect 1880 -2940 1913 -2897
rect 1121 -3011 1154 -2968
rect 1154 -3011 1187 -2968
rect 1088 -3011 1121 -2968
rect 1154 -3011 1187 -2968
rect 1187 -3011 1220 -2968
rect 1220 -3011 1253 -2968
rect 1286 -3011 1319 -2968
rect 1319 -3011 1352 -2968
rect 1352 -3011 1385 -2968
rect 1517 -3011 1550 -2968
rect 1550 -3011 1583 -2968
rect 1484 -3011 1517 -2968
rect 1550 -3011 1583 -2968
rect 1583 -3011 1616 -2968
rect 1616 -3011 1649 -2968
rect 1781 -3011 1814 -2968
rect 1814 -3011 1847 -2968
rect 1748 -3011 1781 -2968
rect 1814 -3011 1847 -2968
rect 1847 -3011 1880 -2968
rect 1880 -3011 1913 -2968
rect 1022 -3082 1055 -3039
rect 1055 -3082 1088 -3039
rect 1088 -3082 1121 -3039
rect 1253 -3082 1286 -3039
rect 1286 -3082 1319 -3039
rect 1220 -3082 1253 -3039
rect 1286 -3082 1319 -3039
rect 1319 -3082 1352 -3039
rect 1352 -3082 1385 -3039
rect 1517 -3082 1550 -3039
rect 1550 -3082 1583 -3039
rect 1484 -3082 1517 -3039
rect 1550 -3082 1583 -3039
rect 1583 -3082 1616 -3039
rect 1616 -3082 1649 -3039
rect 1781 -3082 1814 -3039
rect 1814 -3082 1847 -3039
rect 1748 -3082 1781 -3039
rect 1814 -3082 1847 -3039
rect 1847 -3082 1880 -3039
rect 1880 -3082 1913 -3039
rect 1121 -3153 1154 -3110
rect 1154 -3153 1187 -3110
rect 1088 -3153 1121 -3110
rect 1253 -3153 1286 -3110
rect 1286 -3153 1319 -3110
rect 1220 -3153 1253 -3110
rect 1286 -3153 1319 -3110
rect 1319 -3153 1352 -3110
rect 1352 -3153 1385 -3110
rect 1517 -3153 1550 -3110
rect 1550 -3153 1583 -3110
rect 1484 -3153 1517 -3110
rect 1550 -3153 1583 -3110
rect 1583 -3153 1616 -3110
rect 1616 -3153 1649 -3110
rect 1781 -3153 1814 -3110
rect 1814 -3153 1847 -3110
rect 1748 -3153 1781 -3110
rect 1814 -3153 1847 -3110
rect 1847 -3153 1880 -3110
rect 1880 -3153 1913 -3110
rect 1022 -3224 1055 -3181
rect 1055 -3224 1088 -3181
rect 1088 -3224 1121 -3181
rect 1154 -3224 1187 -3181
rect 1187 -3224 1220 -3181
rect 1220 -3224 1253 -3181
rect 1385 -3224 1418 -3181
rect 1418 -3224 1451 -3181
rect 1352 -3224 1385 -3181
rect 1517 -3224 1550 -3181
rect 1550 -3224 1583 -3181
rect 1484 -3224 1517 -3181
rect 1550 -3224 1583 -3181
rect 1583 -3224 1616 -3181
rect 1616 -3224 1649 -3181
rect 1781 -3224 1814 -3181
rect 1814 -3224 1847 -3181
rect 1748 -3224 1781 -3181
rect 1814 -3224 1847 -3181
rect 1847 -3224 1880 -3181
rect 1880 -3224 1913 -3181
rect 1121 -3295 1154 -3252
rect 1154 -3295 1187 -3252
rect 1088 -3295 1121 -3252
rect 1154 -3295 1187 -3252
rect 1187 -3295 1220 -3252
rect 1220 -3295 1253 -3252
rect 1385 -3295 1418 -3252
rect 1418 -3295 1451 -3252
rect 1352 -3295 1385 -3252
rect 1517 -3295 1550 -3252
rect 1550 -3295 1583 -3252
rect 1484 -3295 1517 -3252
rect 1550 -3295 1583 -3252
rect 1583 -3295 1616 -3252
rect 1616 -3295 1649 -3252
rect 1781 -3295 1814 -3252
rect 1814 -3295 1847 -3252
rect 1748 -3295 1781 -3252
rect 1814 -3295 1847 -3252
rect 1847 -3295 1880 -3252
rect 1880 -3295 1913 -3252
rect 1022 -3366 1055 -3323
rect 1055 -3366 1088 -3323
rect 1088 -3366 1121 -3323
rect 1253 -3366 1286 -3323
rect 1286 -3366 1319 -3323
rect 1220 -3366 1253 -3323
rect 1385 -3366 1418 -3323
rect 1418 -3366 1451 -3323
rect 1352 -3366 1385 -3323
rect 1517 -3366 1550 -3323
rect 1550 -3366 1583 -3323
rect 1484 -3366 1517 -3323
rect 1550 -3366 1583 -3323
rect 1583 -3366 1616 -3323
rect 1616 -3366 1649 -3323
rect 1781 -3366 1814 -3323
rect 1814 -3366 1847 -3323
rect 1748 -3366 1781 -3323
rect 1814 -3366 1847 -3323
rect 1847 -3366 1880 -3323
rect 1880 -3366 1913 -3323
rect 1121 -3437 1154 -3394
rect 1154 -3437 1187 -3394
rect 1088 -3437 1121 -3394
rect 1253 -3437 1286 -3394
rect 1286 -3437 1319 -3394
rect 1220 -3437 1253 -3394
rect 1385 -3437 1418 -3394
rect 1418 -3437 1451 -3394
rect 1352 -3437 1385 -3394
rect 1517 -3437 1550 -3394
rect 1550 -3437 1583 -3394
rect 1484 -3437 1517 -3394
rect 1550 -3437 1583 -3394
rect 1583 -3437 1616 -3394
rect 1616 -3437 1649 -3394
rect 1781 -3437 1814 -3394
rect 1814 -3437 1847 -3394
rect 1748 -3437 1781 -3394
rect 1814 -3437 1847 -3394
rect 1847 -3437 1880 -3394
rect 1880 -3437 1913 -3394
rect 1022 -3508 1055 -3465
rect 1055 -3508 1088 -3465
rect 1088 -3508 1121 -3465
rect 1154 -3508 1187 -3465
rect 1187 -3508 1220 -3465
rect 1220 -3508 1253 -3465
rect 1286 -3508 1319 -3465
rect 1319 -3508 1352 -3465
rect 1352 -3508 1385 -3465
rect 1418 -3508 1451 -3465
rect 1451 -3508 1484 -3465
rect 1484 -3508 1517 -3465
rect 1649 -3508 1682 -3465
rect 1682 -3508 1715 -3465
rect 1616 -3508 1649 -3465
rect 1781 -3508 1814 -3465
rect 1814 -3508 1847 -3465
rect 1748 -3508 1781 -3465
rect 1814 -3508 1847 -3465
rect 1847 -3508 1880 -3465
rect 1880 -3508 1913 -3465
rect 1121 -3579 1154 -3536
rect 1154 -3579 1187 -3536
rect 1088 -3579 1121 -3536
rect 1154 -3579 1187 -3536
rect 1187 -3579 1220 -3536
rect 1220 -3579 1253 -3536
rect 1286 -3579 1319 -3536
rect 1319 -3579 1352 -3536
rect 1352 -3579 1385 -3536
rect 1418 -3579 1451 -3536
rect 1451 -3579 1484 -3536
rect 1484 -3579 1517 -3536
rect 1649 -3579 1682 -3536
rect 1682 -3579 1715 -3536
rect 1616 -3579 1649 -3536
rect 1781 -3579 1814 -3536
rect 1814 -3579 1847 -3536
rect 1748 -3579 1781 -3536
rect 1814 -3579 1847 -3536
rect 1847 -3579 1880 -3536
rect 1880 -3579 1913 -3536
rect 1022 -3650 1055 -3607
rect 1055 -3650 1088 -3607
rect 1088 -3650 1121 -3607
rect 1253 -3650 1286 -3607
rect 1286 -3650 1319 -3607
rect 1220 -3650 1253 -3607
rect 1286 -3650 1319 -3607
rect 1319 -3650 1352 -3607
rect 1352 -3650 1385 -3607
rect 1418 -3650 1451 -3607
rect 1451 -3650 1484 -3607
rect 1484 -3650 1517 -3607
rect 1649 -3650 1682 -3607
rect 1682 -3650 1715 -3607
rect 1616 -3650 1649 -3607
rect 1781 -3650 1814 -3607
rect 1814 -3650 1847 -3607
rect 1748 -3650 1781 -3607
rect 1814 -3650 1847 -3607
rect 1847 -3650 1880 -3607
rect 1880 -3650 1913 -3607
rect 1121 -3721 1154 -3678
rect 1154 -3721 1187 -3678
rect 1088 -3721 1121 -3678
rect 1253 -3721 1286 -3678
rect 1286 -3721 1319 -3678
rect 1220 -3721 1253 -3678
rect 1286 -3721 1319 -3678
rect 1319 -3721 1352 -3678
rect 1352 -3721 1385 -3678
rect 1418 -3721 1451 -3678
rect 1451 -3721 1484 -3678
rect 1484 -3721 1517 -3678
rect 1649 -3721 1682 -3678
rect 1682 -3721 1715 -3678
rect 1616 -3721 1649 -3678
rect 1781 -3721 1814 -3678
rect 1814 -3721 1847 -3678
rect 1748 -3721 1781 -3678
rect 1814 -3721 1847 -3678
rect 1847 -3721 1880 -3678
rect 1880 -3721 1913 -3678
rect 1022 -3792 1055 -3749
rect 1055 -3792 1088 -3749
rect 1088 -3792 1121 -3749
rect 1154 -3792 1187 -3749
rect 1187 -3792 1220 -3749
rect 1220 -3792 1253 -3749
rect 1385 -3792 1418 -3749
rect 1418 -3792 1451 -3749
rect 1352 -3792 1385 -3749
rect 1418 -3792 1451 -3749
rect 1451 -3792 1484 -3749
rect 1484 -3792 1517 -3749
rect 1649 -3792 1682 -3749
rect 1682 -3792 1715 -3749
rect 1616 -3792 1649 -3749
rect 1781 -3792 1814 -3749
rect 1814 -3792 1847 -3749
rect 1748 -3792 1781 -3749
rect 1814 -3792 1847 -3749
rect 1847 -3792 1880 -3749
rect 1880 -3792 1913 -3749
rect 1121 -3863 1154 -3820
rect 1154 -3863 1187 -3820
rect 1088 -3863 1121 -3820
rect 1154 -3863 1187 -3820
rect 1187 -3863 1220 -3820
rect 1220 -3863 1253 -3820
rect 1385 -3863 1418 -3820
rect 1418 -3863 1451 -3820
rect 1352 -3863 1385 -3820
rect 1418 -3863 1451 -3820
rect 1451 -3863 1484 -3820
rect 1484 -3863 1517 -3820
rect 1649 -3863 1682 -3820
rect 1682 -3863 1715 -3820
rect 1616 -3863 1649 -3820
rect 1781 -3863 1814 -3820
rect 1814 -3863 1847 -3820
rect 1748 -3863 1781 -3820
rect 1814 -3863 1847 -3820
rect 1847 -3863 1880 -3820
rect 1880 -3863 1913 -3820
rect 1022 -3934 1055 -3891
rect 1055 -3934 1088 -3891
rect 1088 -3934 1121 -3891
rect 1253 -3934 1286 -3891
rect 1286 -3934 1319 -3891
rect 1220 -3934 1253 -3891
rect 1385 -3934 1418 -3891
rect 1418 -3934 1451 -3891
rect 1352 -3934 1385 -3891
rect 1418 -3934 1451 -3891
rect 1451 -3934 1484 -3891
rect 1484 -3934 1517 -3891
rect 1649 -3934 1682 -3891
rect 1682 -3934 1715 -3891
rect 1616 -3934 1649 -3891
rect 1781 -3934 1814 -3891
rect 1814 -3934 1847 -3891
rect 1748 -3934 1781 -3891
rect 1814 -3934 1847 -3891
rect 1847 -3934 1880 -3891
rect 1880 -3934 1913 -3891
rect 1121 -4005 1154 -3962
rect 1154 -4005 1187 -3962
rect 1088 -4005 1121 -3962
rect 1253 -4005 1286 -3962
rect 1286 -4005 1319 -3962
rect 1220 -4005 1253 -3962
rect 1385 -4005 1418 -3962
rect 1418 -4005 1451 -3962
rect 1352 -4005 1385 -3962
rect 1418 -4005 1451 -3962
rect 1451 -4005 1484 -3962
rect 1484 -4005 1517 -3962
rect 1649 -4005 1682 -3962
rect 1682 -4005 1715 -3962
rect 1616 -4005 1649 -3962
rect 1781 -4005 1814 -3962
rect 1814 -4005 1847 -3962
rect 1748 -4005 1781 -3962
rect 1814 -4005 1847 -3962
rect 1847 -4005 1880 -3962
rect 1880 -4005 1913 -3962
rect 1022 -4076 1055 -4033
rect 1055 -4076 1088 -4033
rect 1088 -4076 1121 -4033
rect 1154 -4076 1187 -4033
rect 1187 -4076 1220 -4033
rect 1220 -4076 1253 -4033
rect 1286 -4076 1319 -4033
rect 1319 -4076 1352 -4033
rect 1352 -4076 1385 -4033
rect 1517 -4076 1550 -4033
rect 1550 -4076 1583 -4033
rect 1484 -4076 1517 -4033
rect 1649 -4076 1682 -4033
rect 1682 -4076 1715 -4033
rect 1616 -4076 1649 -4033
rect 1781 -4076 1814 -4033
rect 1814 -4076 1847 -4033
rect 1748 -4076 1781 -4033
rect 1814 -4076 1847 -4033
rect 1847 -4076 1880 -4033
rect 1880 -4076 1913 -4033
rect 1121 -4147 1154 -4104
rect 1154 -4147 1187 -4104
rect 1088 -4147 1121 -4104
rect 1154 -4147 1187 -4104
rect 1187 -4147 1220 -4104
rect 1220 -4147 1253 -4104
rect 1286 -4147 1319 -4104
rect 1319 -4147 1352 -4104
rect 1352 -4147 1385 -4104
rect 1517 -4147 1550 -4104
rect 1550 -4147 1583 -4104
rect 1484 -4147 1517 -4104
rect 1649 -4147 1682 -4104
rect 1682 -4147 1715 -4104
rect 1616 -4147 1649 -4104
rect 1781 -4147 1814 -4104
rect 1814 -4147 1847 -4104
rect 1748 -4147 1781 -4104
rect 1814 -4147 1847 -4104
rect 1847 -4147 1880 -4104
rect 1880 -4147 1913 -4104
rect 1022 -4218 1055 -4175
rect 1055 -4218 1088 -4175
rect 1088 -4218 1121 -4175
rect 1253 -4218 1286 -4175
rect 1286 -4218 1319 -4175
rect 1220 -4218 1253 -4175
rect 1286 -4218 1319 -4175
rect 1319 -4218 1352 -4175
rect 1352 -4218 1385 -4175
rect 1517 -4218 1550 -4175
rect 1550 -4218 1583 -4175
rect 1484 -4218 1517 -4175
rect 1649 -4218 1682 -4175
rect 1682 -4218 1715 -4175
rect 1616 -4218 1649 -4175
rect 1781 -4218 1814 -4175
rect 1814 -4218 1847 -4175
rect 1748 -4218 1781 -4175
rect 1814 -4218 1847 -4175
rect 1847 -4218 1880 -4175
rect 1880 -4218 1913 -4175
rect 1121 -4289 1154 -4246
rect 1154 -4289 1187 -4246
rect 1088 -4289 1121 -4246
rect 1253 -4289 1286 -4246
rect 1286 -4289 1319 -4246
rect 1220 -4289 1253 -4246
rect 1286 -4289 1319 -4246
rect 1319 -4289 1352 -4246
rect 1352 -4289 1385 -4246
rect 1517 -4289 1550 -4246
rect 1550 -4289 1583 -4246
rect 1484 -4289 1517 -4246
rect 1649 -4289 1682 -4246
rect 1682 -4289 1715 -4246
rect 1616 -4289 1649 -4246
rect 1781 -4289 1814 -4246
rect 1814 -4289 1847 -4246
rect 1748 -4289 1781 -4246
rect 1814 -4289 1847 -4246
rect 1847 -4289 1880 -4246
rect 1880 -4289 1913 -4246
rect 1022 -4360 1055 -4317
rect 1055 -4360 1088 -4317
rect 1088 -4360 1121 -4317
rect 1154 -4360 1187 -4317
rect 1187 -4360 1220 -4317
rect 1220 -4360 1253 -4317
rect 1385 -4360 1418 -4317
rect 1418 -4360 1451 -4317
rect 1352 -4360 1385 -4317
rect 1517 -4360 1550 -4317
rect 1550 -4360 1583 -4317
rect 1484 -4360 1517 -4317
rect 1649 -4360 1682 -4317
rect 1682 -4360 1715 -4317
rect 1616 -4360 1649 -4317
rect 1781 -4360 1814 -4317
rect 1814 -4360 1847 -4317
rect 1748 -4360 1781 -4317
rect 1814 -4360 1847 -4317
rect 1847 -4360 1880 -4317
rect 1880 -4360 1913 -4317
rect 1121 -4431 1154 -4388
rect 1154 -4431 1187 -4388
rect 1088 -4431 1121 -4388
rect 1154 -4431 1187 -4388
rect 1187 -4431 1220 -4388
rect 1220 -4431 1253 -4388
rect 1385 -4431 1418 -4388
rect 1418 -4431 1451 -4388
rect 1352 -4431 1385 -4388
rect 1517 -4431 1550 -4388
rect 1550 -4431 1583 -4388
rect 1484 -4431 1517 -4388
rect 1649 -4431 1682 -4388
rect 1682 -4431 1715 -4388
rect 1616 -4431 1649 -4388
rect 1781 -4431 1814 -4388
rect 1814 -4431 1847 -4388
rect 1748 -4431 1781 -4388
rect 1814 -4431 1847 -4388
rect 1847 -4431 1880 -4388
rect 1880 -4431 1913 -4388
rect 1022 -4502 1055 -4459
rect 1055 -4502 1088 -4459
rect 1088 -4502 1121 -4459
rect 1253 -4502 1286 -4459
rect 1286 -4502 1319 -4459
rect 1220 -4502 1253 -4459
rect 1385 -4502 1418 -4459
rect 1418 -4502 1451 -4459
rect 1352 -4502 1385 -4459
rect 1517 -4502 1550 -4459
rect 1550 -4502 1583 -4459
rect 1484 -4502 1517 -4459
rect 1649 -4502 1682 -4459
rect 1682 -4502 1715 -4459
rect 1616 -4502 1649 -4459
rect 1781 -4502 1814 -4459
rect 1814 -4502 1847 -4459
rect 1748 -4502 1781 -4459
rect 1814 -4502 1847 -4459
rect 1847 -4502 1880 -4459
rect 1880 -4502 1913 -4459
rect 1121 -4573 1154 -4530
rect 1154 -4573 1187 -4530
rect 1088 -4573 1121 -4530
rect 1253 -4573 1286 -4530
rect 1286 -4573 1319 -4530
rect 1220 -4573 1253 -4530
rect 1385 -4573 1418 -4530
rect 1418 -4573 1451 -4530
rect 1352 -4573 1385 -4530
rect 1517 -4573 1550 -4530
rect 1550 -4573 1583 -4530
rect 1484 -4573 1517 -4530
rect 1649 -4573 1682 -4530
rect 1682 -4573 1715 -4530
rect 1616 -4573 1649 -4530
rect 1781 -4573 1814 -4530
rect 1814 -4573 1847 -4530
rect 1748 -4573 1781 -4530
rect 1814 -4573 1847 -4530
rect 1847 -4573 1880 -4530
rect 1880 -4573 1913 -4530
rect 1022 -4644 1055 -4601
rect 1055 -4644 1088 -4601
rect 1088 -4644 1121 -4601
rect 1154 -4644 1187 -4601
rect 1187 -4644 1220 -4601
rect 1220 -4644 1253 -4601
rect 1286 -4644 1319 -4601
rect 1319 -4644 1352 -4601
rect 1352 -4644 1385 -4601
rect 1418 -4644 1451 -4601
rect 1451 -4644 1484 -4601
rect 1484 -4644 1517 -4601
rect 1550 -4644 1583 -4601
rect 1583 -4644 1616 -4601
rect 1616 -4644 1649 -4601
rect 1682 -4644 1715 -4601
rect 1715 -4644 1748 -4601
rect 1748 -4644 1781 -4601
rect 1913 -4644 1946 -4601
rect 1946 -4644 1979 -4601
rect 1880 -4644 1913 -4601
rect 1121 -4715 1154 -4672
rect 1154 -4715 1187 -4672
rect 1088 -4715 1121 -4672
rect 1154 -4715 1187 -4672
rect 1187 -4715 1220 -4672
rect 1220 -4715 1253 -4672
rect 1286 -4715 1319 -4672
rect 1319 -4715 1352 -4672
rect 1352 -4715 1385 -4672
rect 1418 -4715 1451 -4672
rect 1451 -4715 1484 -4672
rect 1484 -4715 1517 -4672
rect 1550 -4715 1583 -4672
rect 1583 -4715 1616 -4672
rect 1616 -4715 1649 -4672
rect 1682 -4715 1715 -4672
rect 1715 -4715 1748 -4672
rect 1748 -4715 1781 -4672
rect 1913 -4715 1946 -4672
rect 1946 -4715 1979 -4672
rect 1880 -4715 1913 -4672
rect 1022 -4786 1055 -4743
rect 1055 -4786 1088 -4743
rect 1088 -4786 1121 -4743
rect 1253 -4786 1286 -4743
rect 1286 -4786 1319 -4743
rect 1220 -4786 1253 -4743
rect 1286 -4786 1319 -4743
rect 1319 -4786 1352 -4743
rect 1352 -4786 1385 -4743
rect 1418 -4786 1451 -4743
rect 1451 -4786 1484 -4743
rect 1484 -4786 1517 -4743
rect 1550 -4786 1583 -4743
rect 1583 -4786 1616 -4743
rect 1616 -4786 1649 -4743
rect 1682 -4786 1715 -4743
rect 1715 -4786 1748 -4743
rect 1748 -4786 1781 -4743
rect 1913 -4786 1946 -4743
rect 1946 -4786 1979 -4743
rect 1880 -4786 1913 -4743
rect 1121 -4857 1154 -4814
rect 1154 -4857 1187 -4814
rect 1088 -4857 1121 -4814
rect 1253 -4857 1286 -4814
rect 1286 -4857 1319 -4814
rect 1220 -4857 1253 -4814
rect 1286 -4857 1319 -4814
rect 1319 -4857 1352 -4814
rect 1352 -4857 1385 -4814
rect 1418 -4857 1451 -4814
rect 1451 -4857 1484 -4814
rect 1484 -4857 1517 -4814
rect 1550 -4857 1583 -4814
rect 1583 -4857 1616 -4814
rect 1616 -4857 1649 -4814
rect 1682 -4857 1715 -4814
rect 1715 -4857 1748 -4814
rect 1748 -4857 1781 -4814
rect 1913 -4857 1946 -4814
rect 1946 -4857 1979 -4814
rect 1880 -4857 1913 -4814
rect 1022 -4928 1055 -4885
rect 1055 -4928 1088 -4885
rect 1088 -4928 1121 -4885
rect 1154 -4928 1187 -4885
rect 1187 -4928 1220 -4885
rect 1220 -4928 1253 -4885
rect 1385 -4928 1418 -4885
rect 1418 -4928 1451 -4885
rect 1352 -4928 1385 -4885
rect 1418 -4928 1451 -4885
rect 1451 -4928 1484 -4885
rect 1484 -4928 1517 -4885
rect 1550 -4928 1583 -4885
rect 1583 -4928 1616 -4885
rect 1616 -4928 1649 -4885
rect 1682 -4928 1715 -4885
rect 1715 -4928 1748 -4885
rect 1748 -4928 1781 -4885
rect 1913 -4928 1946 -4885
rect 1946 -4928 1979 -4885
rect 1880 -4928 1913 -4885
rect 1121 -4999 1154 -4956
rect 1154 -4999 1187 -4956
rect 1088 -4999 1121 -4956
rect 1154 -4999 1187 -4956
rect 1187 -4999 1220 -4956
rect 1220 -4999 1253 -4956
rect 1385 -4999 1418 -4956
rect 1418 -4999 1451 -4956
rect 1352 -4999 1385 -4956
rect 1418 -4999 1451 -4956
rect 1451 -4999 1484 -4956
rect 1484 -4999 1517 -4956
rect 1550 -4999 1583 -4956
rect 1583 -4999 1616 -4956
rect 1616 -4999 1649 -4956
rect 1682 -4999 1715 -4956
rect 1715 -4999 1748 -4956
rect 1748 -4999 1781 -4956
rect 1913 -4999 1946 -4956
rect 1946 -4999 1979 -4956
rect 1880 -4999 1913 -4956
rect 1022 -5070 1055 -5027
rect 1055 -5070 1088 -5027
rect 1088 -5070 1121 -5027
rect 1253 -5070 1286 -5027
rect 1286 -5070 1319 -5027
rect 1220 -5070 1253 -5027
rect 1385 -5070 1418 -5027
rect 1418 -5070 1451 -5027
rect 1352 -5070 1385 -5027
rect 1418 -5070 1451 -5027
rect 1451 -5070 1484 -5027
rect 1484 -5070 1517 -5027
rect 1550 -5070 1583 -5027
rect 1583 -5070 1616 -5027
rect 1616 -5070 1649 -5027
rect 1682 -5070 1715 -5027
rect 1715 -5070 1748 -5027
rect 1748 -5070 1781 -5027
rect 1913 -5070 1946 -5027
rect 1946 -5070 1979 -5027
rect 1880 -5070 1913 -5027
rect 1121 -5141 1154 -5098
rect 1154 -5141 1187 -5098
rect 1088 -5141 1121 -5098
rect 1253 -5141 1286 -5098
rect 1286 -5141 1319 -5098
rect 1220 -5141 1253 -5098
rect 1385 -5141 1418 -5098
rect 1418 -5141 1451 -5098
rect 1352 -5141 1385 -5098
rect 1418 -5141 1451 -5098
rect 1451 -5141 1484 -5098
rect 1484 -5141 1517 -5098
rect 1550 -5141 1583 -5098
rect 1583 -5141 1616 -5098
rect 1616 -5141 1649 -5098
rect 1682 -5141 1715 -5098
rect 1715 -5141 1748 -5098
rect 1748 -5141 1781 -5098
rect 1913 -5141 1946 -5098
rect 1946 -5141 1979 -5098
rect 1880 -5141 1913 -5098
rect 1022 -5212 1055 -5169
rect 1055 -5212 1088 -5169
rect 1088 -5212 1121 -5169
rect 1154 -5212 1187 -5169
rect 1187 -5212 1220 -5169
rect 1220 -5212 1253 -5169
rect 1286 -5212 1319 -5169
rect 1319 -5212 1352 -5169
rect 1352 -5212 1385 -5169
rect 1517 -5212 1550 -5169
rect 1550 -5212 1583 -5169
rect 1484 -5212 1517 -5169
rect 1550 -5212 1583 -5169
rect 1583 -5212 1616 -5169
rect 1616 -5212 1649 -5169
rect 1682 -5212 1715 -5169
rect 1715 -5212 1748 -5169
rect 1748 -5212 1781 -5169
rect 1913 -5212 1946 -5169
rect 1946 -5212 1979 -5169
rect 1880 -5212 1913 -5169
rect 1121 -5283 1154 -5240
rect 1154 -5283 1187 -5240
rect 1088 -5283 1121 -5240
rect 1154 -5283 1187 -5240
rect 1187 -5283 1220 -5240
rect 1220 -5283 1253 -5240
rect 1286 -5283 1319 -5240
rect 1319 -5283 1352 -5240
rect 1352 -5283 1385 -5240
rect 1517 -5283 1550 -5240
rect 1550 -5283 1583 -5240
rect 1484 -5283 1517 -5240
rect 1550 -5283 1583 -5240
rect 1583 -5283 1616 -5240
rect 1616 -5283 1649 -5240
rect 1682 -5283 1715 -5240
rect 1715 -5283 1748 -5240
rect 1748 -5283 1781 -5240
rect 1913 -5283 1946 -5240
rect 1946 -5283 1979 -5240
rect 1880 -5283 1913 -5240
rect 1022 -5354 1055 -5311
rect 1055 -5354 1088 -5311
rect 1088 -5354 1121 -5311
rect 1253 -5354 1286 -5311
rect 1286 -5354 1319 -5311
rect 1220 -5354 1253 -5311
rect 1286 -5354 1319 -5311
rect 1319 -5354 1352 -5311
rect 1352 -5354 1385 -5311
rect 1517 -5354 1550 -5311
rect 1550 -5354 1583 -5311
rect 1484 -5354 1517 -5311
rect 1550 -5354 1583 -5311
rect 1583 -5354 1616 -5311
rect 1616 -5354 1649 -5311
rect 1682 -5354 1715 -5311
rect 1715 -5354 1748 -5311
rect 1748 -5354 1781 -5311
rect 1913 -5354 1946 -5311
rect 1946 -5354 1979 -5311
rect 1880 -5354 1913 -5311
rect 1121 -5425 1154 -5382
rect 1154 -5425 1187 -5382
rect 1088 -5425 1121 -5382
rect 1253 -5425 1286 -5382
rect 1286 -5425 1319 -5382
rect 1220 -5425 1253 -5382
rect 1286 -5425 1319 -5382
rect 1319 -5425 1352 -5382
rect 1352 -5425 1385 -5382
rect 1517 -5425 1550 -5382
rect 1550 -5425 1583 -5382
rect 1484 -5425 1517 -5382
rect 1550 -5425 1583 -5382
rect 1583 -5425 1616 -5382
rect 1616 -5425 1649 -5382
rect 1682 -5425 1715 -5382
rect 1715 -5425 1748 -5382
rect 1748 -5425 1781 -5382
rect 1913 -5425 1946 -5382
rect 1946 -5425 1979 -5382
rect 1880 -5425 1913 -5382
rect 1022 -5496 1055 -5453
rect 1055 -5496 1088 -5453
rect 1088 -5496 1121 -5453
rect 1154 -5496 1187 -5453
rect 1187 -5496 1220 -5453
rect 1220 -5496 1253 -5453
rect 1385 -5496 1418 -5453
rect 1418 -5496 1451 -5453
rect 1352 -5496 1385 -5453
rect 1517 -5496 1550 -5453
rect 1550 -5496 1583 -5453
rect 1484 -5496 1517 -5453
rect 1550 -5496 1583 -5453
rect 1583 -5496 1616 -5453
rect 1616 -5496 1649 -5453
rect 1682 -5496 1715 -5453
rect 1715 -5496 1748 -5453
rect 1748 -5496 1781 -5453
rect 1913 -5496 1946 -5453
rect 1946 -5496 1979 -5453
rect 1880 -5496 1913 -5453
rect 1121 -5567 1154 -5524
rect 1154 -5567 1187 -5524
rect 1088 -5567 1121 -5524
rect 1154 -5567 1187 -5524
rect 1187 -5567 1220 -5524
rect 1220 -5567 1253 -5524
rect 1385 -5567 1418 -5524
rect 1418 -5567 1451 -5524
rect 1352 -5567 1385 -5524
rect 1517 -5567 1550 -5524
rect 1550 -5567 1583 -5524
rect 1484 -5567 1517 -5524
rect 1550 -5567 1583 -5524
rect 1583 -5567 1616 -5524
rect 1616 -5567 1649 -5524
rect 1682 -5567 1715 -5524
rect 1715 -5567 1748 -5524
rect 1748 -5567 1781 -5524
rect 1913 -5567 1946 -5524
rect 1946 -5567 1979 -5524
rect 1880 -5567 1913 -5524
rect 1022 -5638 1055 -5595
rect 1055 -5638 1088 -5595
rect 1088 -5638 1121 -5595
rect 1253 -5638 1286 -5595
rect 1286 -5638 1319 -5595
rect 1220 -5638 1253 -5595
rect 1385 -5638 1418 -5595
rect 1418 -5638 1451 -5595
rect 1352 -5638 1385 -5595
rect 1517 -5638 1550 -5595
rect 1550 -5638 1583 -5595
rect 1484 -5638 1517 -5595
rect 1550 -5638 1583 -5595
rect 1583 -5638 1616 -5595
rect 1616 -5638 1649 -5595
rect 1682 -5638 1715 -5595
rect 1715 -5638 1748 -5595
rect 1748 -5638 1781 -5595
rect 1913 -5638 1946 -5595
rect 1946 -5638 1979 -5595
rect 1880 -5638 1913 -5595
rect 1121 -5709 1154 -5666
rect 1154 -5709 1187 -5666
rect 1088 -5709 1121 -5666
rect 1253 -5709 1286 -5666
rect 1286 -5709 1319 -5666
rect 1220 -5709 1253 -5666
rect 1385 -5709 1418 -5666
rect 1418 -5709 1451 -5666
rect 1352 -5709 1385 -5666
rect 1517 -5709 1550 -5666
rect 1550 -5709 1583 -5666
rect 1484 -5709 1517 -5666
rect 1550 -5709 1583 -5666
rect 1583 -5709 1616 -5666
rect 1616 -5709 1649 -5666
rect 1682 -5709 1715 -5666
rect 1715 -5709 1748 -5666
rect 1748 -5709 1781 -5666
rect 1913 -5709 1946 -5666
rect 1946 -5709 1979 -5666
rect 1880 -5709 1913 -5666
rect 1022 -5780 1055 -5737
rect 1055 -5780 1088 -5737
rect 1088 -5780 1121 -5737
rect 1154 -5780 1187 -5737
rect 1187 -5780 1220 -5737
rect 1220 -5780 1253 -5737
rect 1286 -5780 1319 -5737
rect 1319 -5780 1352 -5737
rect 1352 -5780 1385 -5737
rect 1418 -5780 1451 -5737
rect 1451 -5780 1484 -5737
rect 1484 -5780 1517 -5737
rect 1649 -5780 1682 -5737
rect 1682 -5780 1715 -5737
rect 1616 -5780 1649 -5737
rect 1682 -5780 1715 -5737
rect 1715 -5780 1748 -5737
rect 1748 -5780 1781 -5737
rect 1913 -5780 1946 -5737
rect 1946 -5780 1979 -5737
rect 1880 -5780 1913 -5737
rect 1121 -5851 1154 -5808
rect 1154 -5851 1187 -5808
rect 1088 -5851 1121 -5808
rect 1154 -5851 1187 -5808
rect 1187 -5851 1220 -5808
rect 1220 -5851 1253 -5808
rect 1286 -5851 1319 -5808
rect 1319 -5851 1352 -5808
rect 1352 -5851 1385 -5808
rect 1418 -5851 1451 -5808
rect 1451 -5851 1484 -5808
rect 1484 -5851 1517 -5808
rect 1649 -5851 1682 -5808
rect 1682 -5851 1715 -5808
rect 1616 -5851 1649 -5808
rect 1682 -5851 1715 -5808
rect 1715 -5851 1748 -5808
rect 1748 -5851 1781 -5808
rect 1913 -5851 1946 -5808
rect 1946 -5851 1979 -5808
rect 1880 -5851 1913 -5808
rect 1022 -5922 1055 -5879
rect 1055 -5922 1088 -5879
rect 1088 -5922 1121 -5879
rect 1253 -5922 1286 -5879
rect 1286 -5922 1319 -5879
rect 1220 -5922 1253 -5879
rect 1286 -5922 1319 -5879
rect 1319 -5922 1352 -5879
rect 1352 -5922 1385 -5879
rect 1418 -5922 1451 -5879
rect 1451 -5922 1484 -5879
rect 1484 -5922 1517 -5879
rect 1649 -5922 1682 -5879
rect 1682 -5922 1715 -5879
rect 1616 -5922 1649 -5879
rect 1682 -5922 1715 -5879
rect 1715 -5922 1748 -5879
rect 1748 -5922 1781 -5879
rect 1913 -5922 1946 -5879
rect 1946 -5922 1979 -5879
rect 1880 -5922 1913 -5879
rect 1121 -5993 1154 -5950
rect 1154 -5993 1187 -5950
rect 1088 -5993 1121 -5950
rect 1253 -5993 1286 -5950
rect 1286 -5993 1319 -5950
rect 1220 -5993 1253 -5950
rect 1286 -5993 1319 -5950
rect 1319 -5993 1352 -5950
rect 1352 -5993 1385 -5950
rect 1418 -5993 1451 -5950
rect 1451 -5993 1484 -5950
rect 1484 -5993 1517 -5950
rect 1649 -5993 1682 -5950
rect 1682 -5993 1715 -5950
rect 1616 -5993 1649 -5950
rect 1682 -5993 1715 -5950
rect 1715 -5993 1748 -5950
rect 1748 -5993 1781 -5950
rect 1913 -5993 1946 -5950
rect 1946 -5993 1979 -5950
rect 1880 -5993 1913 -5950
rect 1022 -6064 1055 -6021
rect 1055 -6064 1088 -6021
rect 1088 -6064 1121 -6021
rect 1154 -6064 1187 -6021
rect 1187 -6064 1220 -6021
rect 1220 -6064 1253 -6021
rect 1385 -6064 1418 -6021
rect 1418 -6064 1451 -6021
rect 1352 -6064 1385 -6021
rect 1418 -6064 1451 -6021
rect 1451 -6064 1484 -6021
rect 1484 -6064 1517 -6021
rect 1649 -6064 1682 -6021
rect 1682 -6064 1715 -6021
rect 1616 -6064 1649 -6021
rect 1682 -6064 1715 -6021
rect 1715 -6064 1748 -6021
rect 1748 -6064 1781 -6021
rect 1913 -6064 1946 -6021
rect 1946 -6064 1979 -6021
rect 1880 -6064 1913 -6021
rect 1121 -6135 1154 -6092
rect 1154 -6135 1187 -6092
rect 1088 -6135 1121 -6092
rect 1154 -6135 1187 -6092
rect 1187 -6135 1220 -6092
rect 1220 -6135 1253 -6092
rect 1385 -6135 1418 -6092
rect 1418 -6135 1451 -6092
rect 1352 -6135 1385 -6092
rect 1418 -6135 1451 -6092
rect 1451 -6135 1484 -6092
rect 1484 -6135 1517 -6092
rect 1649 -6135 1682 -6092
rect 1682 -6135 1715 -6092
rect 1616 -6135 1649 -6092
rect 1682 -6135 1715 -6092
rect 1715 -6135 1748 -6092
rect 1748 -6135 1781 -6092
rect 1913 -6135 1946 -6092
rect 1946 -6135 1979 -6092
rect 1880 -6135 1913 -6092
rect 1022 -6206 1055 -6163
rect 1055 -6206 1088 -6163
rect 1088 -6206 1121 -6163
rect 1253 -6206 1286 -6163
rect 1286 -6206 1319 -6163
rect 1220 -6206 1253 -6163
rect 1385 -6206 1418 -6163
rect 1418 -6206 1451 -6163
rect 1352 -6206 1385 -6163
rect 1418 -6206 1451 -6163
rect 1451 -6206 1484 -6163
rect 1484 -6206 1517 -6163
rect 1649 -6206 1682 -6163
rect 1682 -6206 1715 -6163
rect 1616 -6206 1649 -6163
rect 1682 -6206 1715 -6163
rect 1715 -6206 1748 -6163
rect 1748 -6206 1781 -6163
rect 1913 -6206 1946 -6163
rect 1946 -6206 1979 -6163
rect 1880 -6206 1913 -6163
rect 1121 -6277 1154 -6234
rect 1154 -6277 1187 -6234
rect 1088 -6277 1121 -6234
rect 1253 -6277 1286 -6234
rect 1286 -6277 1319 -6234
rect 1220 -6277 1253 -6234
rect 1385 -6277 1418 -6234
rect 1418 -6277 1451 -6234
rect 1352 -6277 1385 -6234
rect 1418 -6277 1451 -6234
rect 1451 -6277 1484 -6234
rect 1484 -6277 1517 -6234
rect 1649 -6277 1682 -6234
rect 1682 -6277 1715 -6234
rect 1616 -6277 1649 -6234
rect 1682 -6277 1715 -6234
rect 1715 -6277 1748 -6234
rect 1748 -6277 1781 -6234
rect 1913 -6277 1946 -6234
rect 1946 -6277 1979 -6234
rect 1880 -6277 1913 -6234
rect 1022 -6348 1055 -6305
rect 1055 -6348 1088 -6305
rect 1088 -6348 1121 -6305
rect 1154 -6348 1187 -6305
rect 1187 -6348 1220 -6305
rect 1220 -6348 1253 -6305
rect 1286 -6348 1319 -6305
rect 1319 -6348 1352 -6305
rect 1352 -6348 1385 -6305
rect 1517 -6348 1550 -6305
rect 1550 -6348 1583 -6305
rect 1484 -6348 1517 -6305
rect 1649 -6348 1682 -6305
rect 1682 -6348 1715 -6305
rect 1616 -6348 1649 -6305
rect 1682 -6348 1715 -6305
rect 1715 -6348 1748 -6305
rect 1748 -6348 1781 -6305
rect 1913 -6348 1946 -6305
rect 1946 -6348 1979 -6305
rect 1880 -6348 1913 -6305
rect 1121 -6419 1154 -6376
rect 1154 -6419 1187 -6376
rect 1088 -6419 1121 -6376
rect 1154 -6419 1187 -6376
rect 1187 -6419 1220 -6376
rect 1220 -6419 1253 -6376
rect 1286 -6419 1319 -6376
rect 1319 -6419 1352 -6376
rect 1352 -6419 1385 -6376
rect 1517 -6419 1550 -6376
rect 1550 -6419 1583 -6376
rect 1484 -6419 1517 -6376
rect 1649 -6419 1682 -6376
rect 1682 -6419 1715 -6376
rect 1616 -6419 1649 -6376
rect 1682 -6419 1715 -6376
rect 1715 -6419 1748 -6376
rect 1748 -6419 1781 -6376
rect 1913 -6419 1946 -6376
rect 1946 -6419 1979 -6376
rect 1880 -6419 1913 -6376
rect 1022 -6490 1055 -6447
rect 1055 -6490 1088 -6447
rect 1088 -6490 1121 -6447
rect 1253 -6490 1286 -6447
rect 1286 -6490 1319 -6447
rect 1220 -6490 1253 -6447
rect 1286 -6490 1319 -6447
rect 1319 -6490 1352 -6447
rect 1352 -6490 1385 -6447
rect 1517 -6490 1550 -6447
rect 1550 -6490 1583 -6447
rect 1484 -6490 1517 -6447
rect 1649 -6490 1682 -6447
rect 1682 -6490 1715 -6447
rect 1616 -6490 1649 -6447
rect 1682 -6490 1715 -6447
rect 1715 -6490 1748 -6447
rect 1748 -6490 1781 -6447
rect 1913 -6490 1946 -6447
rect 1946 -6490 1979 -6447
rect 1880 -6490 1913 -6447
rect 1121 -6561 1154 -6518
rect 1154 -6561 1187 -6518
rect 1088 -6561 1121 -6518
rect 1253 -6561 1286 -6518
rect 1286 -6561 1319 -6518
rect 1220 -6561 1253 -6518
rect 1286 -6561 1319 -6518
rect 1319 -6561 1352 -6518
rect 1352 -6561 1385 -6518
rect 1517 -6561 1550 -6518
rect 1550 -6561 1583 -6518
rect 1484 -6561 1517 -6518
rect 1649 -6561 1682 -6518
rect 1682 -6561 1715 -6518
rect 1616 -6561 1649 -6518
rect 1682 -6561 1715 -6518
rect 1715 -6561 1748 -6518
rect 1748 -6561 1781 -6518
rect 1913 -6561 1946 -6518
rect 1946 -6561 1979 -6518
rect 1880 -6561 1913 -6518
rect 1022 -6632 1055 -6589
rect 1055 -6632 1088 -6589
rect 1088 -6632 1121 -6589
rect 1154 -6632 1187 -6589
rect 1187 -6632 1220 -6589
rect 1220 -6632 1253 -6589
rect 1385 -6632 1418 -6589
rect 1418 -6632 1451 -6589
rect 1352 -6632 1385 -6589
rect 1517 -6632 1550 -6589
rect 1550 -6632 1583 -6589
rect 1484 -6632 1517 -6589
rect 1649 -6632 1682 -6589
rect 1682 -6632 1715 -6589
rect 1616 -6632 1649 -6589
rect 1682 -6632 1715 -6589
rect 1715 -6632 1748 -6589
rect 1748 -6632 1781 -6589
rect 1913 -6632 1946 -6589
rect 1946 -6632 1979 -6589
rect 1880 -6632 1913 -6589
rect 1121 -6703 1154 -6660
rect 1154 -6703 1187 -6660
rect 1088 -6703 1121 -6660
rect 1154 -6703 1187 -6660
rect 1187 -6703 1220 -6660
rect 1220 -6703 1253 -6660
rect 1385 -6703 1418 -6660
rect 1418 -6703 1451 -6660
rect 1352 -6703 1385 -6660
rect 1517 -6703 1550 -6660
rect 1550 -6703 1583 -6660
rect 1484 -6703 1517 -6660
rect 1649 -6703 1682 -6660
rect 1682 -6703 1715 -6660
rect 1616 -6703 1649 -6660
rect 1682 -6703 1715 -6660
rect 1715 -6703 1748 -6660
rect 1748 -6703 1781 -6660
rect 1913 -6703 1946 -6660
rect 1946 -6703 1979 -6660
rect 1880 -6703 1913 -6660
rect 1022 -6774 1055 -6731
rect 1055 -6774 1088 -6731
rect 1088 -6774 1121 -6731
rect 1253 -6774 1286 -6731
rect 1286 -6774 1319 -6731
rect 1220 -6774 1253 -6731
rect 1385 -6774 1418 -6731
rect 1418 -6774 1451 -6731
rect 1352 -6774 1385 -6731
rect 1517 -6774 1550 -6731
rect 1550 -6774 1583 -6731
rect 1484 -6774 1517 -6731
rect 1649 -6774 1682 -6731
rect 1682 -6774 1715 -6731
rect 1616 -6774 1649 -6731
rect 1682 -6774 1715 -6731
rect 1715 -6774 1748 -6731
rect 1748 -6774 1781 -6731
rect 1913 -6774 1946 -6731
rect 1946 -6774 1979 -6731
rect 1880 -6774 1913 -6731
rect 1121 -6845 1154 -6802
rect 1154 -6845 1187 -6802
rect 1088 -6845 1121 -6802
rect 1253 -6845 1286 -6802
rect 1286 -6845 1319 -6802
rect 1220 -6845 1253 -6802
rect 1385 -6845 1418 -6802
rect 1418 -6845 1451 -6802
rect 1352 -6845 1385 -6802
rect 1517 -6845 1550 -6802
rect 1550 -6845 1583 -6802
rect 1484 -6845 1517 -6802
rect 1649 -6845 1682 -6802
rect 1682 -6845 1715 -6802
rect 1616 -6845 1649 -6802
rect 1682 -6845 1715 -6802
rect 1715 -6845 1748 -6802
rect 1748 -6845 1781 -6802
rect 1913 -6845 1946 -6802
rect 1946 -6845 1979 -6802
rect 1880 -6845 1913 -6802
rect 1022 -6916 1055 -6873
rect 1055 -6916 1088 -6873
rect 1088 -6916 1121 -6873
rect 1154 -6916 1187 -6873
rect 1187 -6916 1220 -6873
rect 1220 -6916 1253 -6873
rect 1286 -6916 1319 -6873
rect 1319 -6916 1352 -6873
rect 1352 -6916 1385 -6873
rect 1418 -6916 1451 -6873
rect 1451 -6916 1484 -6873
rect 1484 -6916 1517 -6873
rect 1550 -6916 1583 -6873
rect 1583 -6916 1616 -6873
rect 1616 -6916 1649 -6873
rect 1781 -6916 1814 -6873
rect 1814 -6916 1847 -6873
rect 1748 -6916 1781 -6873
rect 1913 -6916 1946 -6873
rect 1946 -6916 1979 -6873
rect 1880 -6916 1913 -6873
rect 1121 -6987 1154 -6944
rect 1154 -6987 1187 -6944
rect 1088 -6987 1121 -6944
rect 1154 -6987 1187 -6944
rect 1187 -6987 1220 -6944
rect 1220 -6987 1253 -6944
rect 1286 -6987 1319 -6944
rect 1319 -6987 1352 -6944
rect 1352 -6987 1385 -6944
rect 1418 -6987 1451 -6944
rect 1451 -6987 1484 -6944
rect 1484 -6987 1517 -6944
rect 1550 -6987 1583 -6944
rect 1583 -6987 1616 -6944
rect 1616 -6987 1649 -6944
rect 1781 -6987 1814 -6944
rect 1814 -6987 1847 -6944
rect 1748 -6987 1781 -6944
rect 1913 -6987 1946 -6944
rect 1946 -6987 1979 -6944
rect 1880 -6987 1913 -6944
rect 1022 -7058 1055 -7015
rect 1055 -7058 1088 -7015
rect 1088 -7058 1121 -7015
rect 1253 -7058 1286 -7015
rect 1286 -7058 1319 -7015
rect 1220 -7058 1253 -7015
rect 1286 -7058 1319 -7015
rect 1319 -7058 1352 -7015
rect 1352 -7058 1385 -7015
rect 1418 -7058 1451 -7015
rect 1451 -7058 1484 -7015
rect 1484 -7058 1517 -7015
rect 1550 -7058 1583 -7015
rect 1583 -7058 1616 -7015
rect 1616 -7058 1649 -7015
rect 1781 -7058 1814 -7015
rect 1814 -7058 1847 -7015
rect 1748 -7058 1781 -7015
rect 1913 -7058 1946 -7015
rect 1946 -7058 1979 -7015
rect 1880 -7058 1913 -7015
rect 1121 -7129 1154 -7086
rect 1154 -7129 1187 -7086
rect 1088 -7129 1121 -7086
rect 1253 -7129 1286 -7086
rect 1286 -7129 1319 -7086
rect 1220 -7129 1253 -7086
rect 1286 -7129 1319 -7086
rect 1319 -7129 1352 -7086
rect 1352 -7129 1385 -7086
rect 1418 -7129 1451 -7086
rect 1451 -7129 1484 -7086
rect 1484 -7129 1517 -7086
rect 1550 -7129 1583 -7086
rect 1583 -7129 1616 -7086
rect 1616 -7129 1649 -7086
rect 1781 -7129 1814 -7086
rect 1814 -7129 1847 -7086
rect 1748 -7129 1781 -7086
rect 1913 -7129 1946 -7086
rect 1946 -7129 1979 -7086
rect 1880 -7129 1913 -7086
rect 1022 -7200 1055 -7157
rect 1055 -7200 1088 -7157
rect 1088 -7200 1121 -7157
rect 1154 -7200 1187 -7157
rect 1187 -7200 1220 -7157
rect 1220 -7200 1253 -7157
rect 1385 -7200 1418 -7157
rect 1418 -7200 1451 -7157
rect 1352 -7200 1385 -7157
rect 1418 -7200 1451 -7157
rect 1451 -7200 1484 -7157
rect 1484 -7200 1517 -7157
rect 1550 -7200 1583 -7157
rect 1583 -7200 1616 -7157
rect 1616 -7200 1649 -7157
rect 1781 -7200 1814 -7157
rect 1814 -7200 1847 -7157
rect 1748 -7200 1781 -7157
rect 1913 -7200 1946 -7157
rect 1946 -7200 1979 -7157
rect 1880 -7200 1913 -7157
rect 1121 -7271 1154 -7228
rect 1154 -7271 1187 -7228
rect 1088 -7271 1121 -7228
rect 1154 -7271 1187 -7228
rect 1187 -7271 1220 -7228
rect 1220 -7271 1253 -7228
rect 1385 -7271 1418 -7228
rect 1418 -7271 1451 -7228
rect 1352 -7271 1385 -7228
rect 1418 -7271 1451 -7228
rect 1451 -7271 1484 -7228
rect 1484 -7271 1517 -7228
rect 1550 -7271 1583 -7228
rect 1583 -7271 1616 -7228
rect 1616 -7271 1649 -7228
rect 1781 -7271 1814 -7228
rect 1814 -7271 1847 -7228
rect 1748 -7271 1781 -7228
rect 1913 -7271 1946 -7228
rect 1946 -7271 1979 -7228
rect 1880 -7271 1913 -7228
rect 1022 -7342 1055 -7299
rect 1055 -7342 1088 -7299
rect 1088 -7342 1121 -7299
rect 1253 -7342 1286 -7299
rect 1286 -7342 1319 -7299
rect 1220 -7342 1253 -7299
rect 1385 -7342 1418 -7299
rect 1418 -7342 1451 -7299
rect 1352 -7342 1385 -7299
rect 1418 -7342 1451 -7299
rect 1451 -7342 1484 -7299
rect 1484 -7342 1517 -7299
rect 1550 -7342 1583 -7299
rect 1583 -7342 1616 -7299
rect 1616 -7342 1649 -7299
rect 1781 -7342 1814 -7299
rect 1814 -7342 1847 -7299
rect 1748 -7342 1781 -7299
rect 1913 -7342 1946 -7299
rect 1946 -7342 1979 -7299
rect 1880 -7342 1913 -7299
rect 1121 -7413 1154 -7370
rect 1154 -7413 1187 -7370
rect 1088 -7413 1121 -7370
rect 1253 -7413 1286 -7370
rect 1286 -7413 1319 -7370
rect 1220 -7413 1253 -7370
rect 1385 -7413 1418 -7370
rect 1418 -7413 1451 -7370
rect 1352 -7413 1385 -7370
rect 1418 -7413 1451 -7370
rect 1451 -7413 1484 -7370
rect 1484 -7413 1517 -7370
rect 1550 -7413 1583 -7370
rect 1583 -7413 1616 -7370
rect 1616 -7413 1649 -7370
rect 1781 -7413 1814 -7370
rect 1814 -7413 1847 -7370
rect 1748 -7413 1781 -7370
rect 1913 -7413 1946 -7370
rect 1946 -7413 1979 -7370
rect 1880 -7413 1913 -7370
rect 1022 -7484 1055 -7441
rect 1055 -7484 1088 -7441
rect 1088 -7484 1121 -7441
rect 1154 -7484 1187 -7441
rect 1187 -7484 1220 -7441
rect 1220 -7484 1253 -7441
rect 1286 -7484 1319 -7441
rect 1319 -7484 1352 -7441
rect 1352 -7484 1385 -7441
rect 1517 -7484 1550 -7441
rect 1550 -7484 1583 -7441
rect 1484 -7484 1517 -7441
rect 1550 -7484 1583 -7441
rect 1583 -7484 1616 -7441
rect 1616 -7484 1649 -7441
rect 1781 -7484 1814 -7441
rect 1814 -7484 1847 -7441
rect 1748 -7484 1781 -7441
rect 1913 -7484 1946 -7441
rect 1946 -7484 1979 -7441
rect 1880 -7484 1913 -7441
rect 1121 -7555 1154 -7512
rect 1154 -7555 1187 -7512
rect 1088 -7555 1121 -7512
rect 1154 -7555 1187 -7512
rect 1187 -7555 1220 -7512
rect 1220 -7555 1253 -7512
rect 1286 -7555 1319 -7512
rect 1319 -7555 1352 -7512
rect 1352 -7555 1385 -7512
rect 1517 -7555 1550 -7512
rect 1550 -7555 1583 -7512
rect 1484 -7555 1517 -7512
rect 1550 -7555 1583 -7512
rect 1583 -7555 1616 -7512
rect 1616 -7555 1649 -7512
rect 1781 -7555 1814 -7512
rect 1814 -7555 1847 -7512
rect 1748 -7555 1781 -7512
rect 1913 -7555 1946 -7512
rect 1946 -7555 1979 -7512
rect 1880 -7555 1913 -7512
rect 1022 -7626 1055 -7583
rect 1055 -7626 1088 -7583
rect 1088 -7626 1121 -7583
rect 1253 -7626 1286 -7583
rect 1286 -7626 1319 -7583
rect 1220 -7626 1253 -7583
rect 1286 -7626 1319 -7583
rect 1319 -7626 1352 -7583
rect 1352 -7626 1385 -7583
rect 1517 -7626 1550 -7583
rect 1550 -7626 1583 -7583
rect 1484 -7626 1517 -7583
rect 1550 -7626 1583 -7583
rect 1583 -7626 1616 -7583
rect 1616 -7626 1649 -7583
rect 1781 -7626 1814 -7583
rect 1814 -7626 1847 -7583
rect 1748 -7626 1781 -7583
rect 1913 -7626 1946 -7583
rect 1946 -7626 1979 -7583
rect 1880 -7626 1913 -7583
rect 1121 -7697 1154 -7654
rect 1154 -7697 1187 -7654
rect 1088 -7697 1121 -7654
rect 1253 -7697 1286 -7654
rect 1286 -7697 1319 -7654
rect 1220 -7697 1253 -7654
rect 1286 -7697 1319 -7654
rect 1319 -7697 1352 -7654
rect 1352 -7697 1385 -7654
rect 1517 -7697 1550 -7654
rect 1550 -7697 1583 -7654
rect 1484 -7697 1517 -7654
rect 1550 -7697 1583 -7654
rect 1583 -7697 1616 -7654
rect 1616 -7697 1649 -7654
rect 1781 -7697 1814 -7654
rect 1814 -7697 1847 -7654
rect 1748 -7697 1781 -7654
rect 1913 -7697 1946 -7654
rect 1946 -7697 1979 -7654
rect 1880 -7697 1913 -7654
rect 1022 -7768 1055 -7725
rect 1055 -7768 1088 -7725
rect 1088 -7768 1121 -7725
rect 1154 -7768 1187 -7725
rect 1187 -7768 1220 -7725
rect 1220 -7768 1253 -7725
rect 1385 -7768 1418 -7725
rect 1418 -7768 1451 -7725
rect 1352 -7768 1385 -7725
rect 1517 -7768 1550 -7725
rect 1550 -7768 1583 -7725
rect 1484 -7768 1517 -7725
rect 1550 -7768 1583 -7725
rect 1583 -7768 1616 -7725
rect 1616 -7768 1649 -7725
rect 1781 -7768 1814 -7725
rect 1814 -7768 1847 -7725
rect 1748 -7768 1781 -7725
rect 1913 -7768 1946 -7725
rect 1946 -7768 1979 -7725
rect 1880 -7768 1913 -7725
rect 1121 -7839 1154 -7796
rect 1154 -7839 1187 -7796
rect 1088 -7839 1121 -7796
rect 1154 -7839 1187 -7796
rect 1187 -7839 1220 -7796
rect 1220 -7839 1253 -7796
rect 1385 -7839 1418 -7796
rect 1418 -7839 1451 -7796
rect 1352 -7839 1385 -7796
rect 1517 -7839 1550 -7796
rect 1550 -7839 1583 -7796
rect 1484 -7839 1517 -7796
rect 1550 -7839 1583 -7796
rect 1583 -7839 1616 -7796
rect 1616 -7839 1649 -7796
rect 1781 -7839 1814 -7796
rect 1814 -7839 1847 -7796
rect 1748 -7839 1781 -7796
rect 1913 -7839 1946 -7796
rect 1946 -7839 1979 -7796
rect 1880 -7839 1913 -7796
rect 1022 -7910 1055 -7867
rect 1055 -7910 1088 -7867
rect 1088 -7910 1121 -7867
rect 1253 -7910 1286 -7867
rect 1286 -7910 1319 -7867
rect 1220 -7910 1253 -7867
rect 1385 -7910 1418 -7867
rect 1418 -7910 1451 -7867
rect 1352 -7910 1385 -7867
rect 1517 -7910 1550 -7867
rect 1550 -7910 1583 -7867
rect 1484 -7910 1517 -7867
rect 1550 -7910 1583 -7867
rect 1583 -7910 1616 -7867
rect 1616 -7910 1649 -7867
rect 1781 -7910 1814 -7867
rect 1814 -7910 1847 -7867
rect 1748 -7910 1781 -7867
rect 1913 -7910 1946 -7867
rect 1946 -7910 1979 -7867
rect 1880 -7910 1913 -7867
rect 1121 -7981 1154 -7938
rect 1154 -7981 1187 -7938
rect 1088 -7981 1121 -7938
rect 1253 -7981 1286 -7938
rect 1286 -7981 1319 -7938
rect 1220 -7981 1253 -7938
rect 1385 -7981 1418 -7938
rect 1418 -7981 1451 -7938
rect 1352 -7981 1385 -7938
rect 1517 -7981 1550 -7938
rect 1550 -7981 1583 -7938
rect 1484 -7981 1517 -7938
rect 1550 -7981 1583 -7938
rect 1583 -7981 1616 -7938
rect 1616 -7981 1649 -7938
rect 1781 -7981 1814 -7938
rect 1814 -7981 1847 -7938
rect 1748 -7981 1781 -7938
rect 1913 -7981 1946 -7938
rect 1946 -7981 1979 -7938
rect 1880 -7981 1913 -7938
rect 1022 -8052 1055 -8009
rect 1055 -8052 1088 -8009
rect 1088 -8052 1121 -8009
rect 1154 -8052 1187 -8009
rect 1187 -8052 1220 -8009
rect 1220 -8052 1253 -8009
rect 1286 -8052 1319 -8009
rect 1319 -8052 1352 -8009
rect 1352 -8052 1385 -8009
rect 1418 -8052 1451 -8009
rect 1451 -8052 1484 -8009
rect 1484 -8052 1517 -8009
rect 1649 -8052 1682 -8009
rect 1682 -8052 1715 -8009
rect 1616 -8052 1649 -8009
rect 1781 -8052 1814 -8009
rect 1814 -8052 1847 -8009
rect 1748 -8052 1781 -8009
rect 1913 -8052 1946 -8009
rect 1946 -8052 1979 -8009
rect 1880 -8052 1913 -8009
rect 1121 -8123 1154 -8080
rect 1154 -8123 1187 -8080
rect 1088 -8123 1121 -8080
rect 1154 -8123 1187 -8080
rect 1187 -8123 1220 -8080
rect 1220 -8123 1253 -8080
rect 1286 -8123 1319 -8080
rect 1319 -8123 1352 -8080
rect 1352 -8123 1385 -8080
rect 1418 -8123 1451 -8080
rect 1451 -8123 1484 -8080
rect 1484 -8123 1517 -8080
rect 1649 -8123 1682 -8080
rect 1682 -8123 1715 -8080
rect 1616 -8123 1649 -8080
rect 1781 -8123 1814 -8080
rect 1814 -8123 1847 -8080
rect 1748 -8123 1781 -8080
rect 1913 -8123 1946 -8080
rect 1946 -8123 1979 -8080
rect 1880 -8123 1913 -8080
rect 1022 -8194 1055 -8151
rect 1055 -8194 1088 -8151
rect 1088 -8194 1121 -8151
rect 1253 -8194 1286 -8151
rect 1286 -8194 1319 -8151
rect 1220 -8194 1253 -8151
rect 1286 -8194 1319 -8151
rect 1319 -8194 1352 -8151
rect 1352 -8194 1385 -8151
rect 1418 -8194 1451 -8151
rect 1451 -8194 1484 -8151
rect 1484 -8194 1517 -8151
rect 1649 -8194 1682 -8151
rect 1682 -8194 1715 -8151
rect 1616 -8194 1649 -8151
rect 1781 -8194 1814 -8151
rect 1814 -8194 1847 -8151
rect 1748 -8194 1781 -8151
rect 1913 -8194 1946 -8151
rect 1946 -8194 1979 -8151
rect 1880 -8194 1913 -8151
rect 1121 -8265 1154 -8222
rect 1154 -8265 1187 -8222
rect 1088 -8265 1121 -8222
rect 1253 -8265 1286 -8222
rect 1286 -8265 1319 -8222
rect 1220 -8265 1253 -8222
rect 1286 -8265 1319 -8222
rect 1319 -8265 1352 -8222
rect 1352 -8265 1385 -8222
rect 1418 -8265 1451 -8222
rect 1451 -8265 1484 -8222
rect 1484 -8265 1517 -8222
rect 1649 -8265 1682 -8222
rect 1682 -8265 1715 -8222
rect 1616 -8265 1649 -8222
rect 1781 -8265 1814 -8222
rect 1814 -8265 1847 -8222
rect 1748 -8265 1781 -8222
rect 1913 -8265 1946 -8222
rect 1946 -8265 1979 -8222
rect 1880 -8265 1913 -8222
rect 1022 -8336 1055 -8293
rect 1055 -8336 1088 -8293
rect 1088 -8336 1121 -8293
rect 1154 -8336 1187 -8293
rect 1187 -8336 1220 -8293
rect 1220 -8336 1253 -8293
rect 1385 -8336 1418 -8293
rect 1418 -8336 1451 -8293
rect 1352 -8336 1385 -8293
rect 1418 -8336 1451 -8293
rect 1451 -8336 1484 -8293
rect 1484 -8336 1517 -8293
rect 1649 -8336 1682 -8293
rect 1682 -8336 1715 -8293
rect 1616 -8336 1649 -8293
rect 1781 -8336 1814 -8293
rect 1814 -8336 1847 -8293
rect 1748 -8336 1781 -8293
rect 1913 -8336 1946 -8293
rect 1946 -8336 1979 -8293
rect 1880 -8336 1913 -8293
rect 1121 -8407 1154 -8364
rect 1154 -8407 1187 -8364
rect 1088 -8407 1121 -8364
rect 1154 -8407 1187 -8364
rect 1187 -8407 1220 -8364
rect 1220 -8407 1253 -8364
rect 1385 -8407 1418 -8364
rect 1418 -8407 1451 -8364
rect 1352 -8407 1385 -8364
rect 1418 -8407 1451 -8364
rect 1451 -8407 1484 -8364
rect 1484 -8407 1517 -8364
rect 1649 -8407 1682 -8364
rect 1682 -8407 1715 -8364
rect 1616 -8407 1649 -8364
rect 1781 -8407 1814 -8364
rect 1814 -8407 1847 -8364
rect 1748 -8407 1781 -8364
rect 1913 -8407 1946 -8364
rect 1946 -8407 1979 -8364
rect 1880 -8407 1913 -8364
rect 1022 -8478 1055 -8435
rect 1055 -8478 1088 -8435
rect 1088 -8478 1121 -8435
rect 1253 -8478 1286 -8435
rect 1286 -8478 1319 -8435
rect 1220 -8478 1253 -8435
rect 1385 -8478 1418 -8435
rect 1418 -8478 1451 -8435
rect 1352 -8478 1385 -8435
rect 1418 -8478 1451 -8435
rect 1451 -8478 1484 -8435
rect 1484 -8478 1517 -8435
rect 1649 -8478 1682 -8435
rect 1682 -8478 1715 -8435
rect 1616 -8478 1649 -8435
rect 1781 -8478 1814 -8435
rect 1814 -8478 1847 -8435
rect 1748 -8478 1781 -8435
rect 1913 -8478 1946 -8435
rect 1946 -8478 1979 -8435
rect 1880 -8478 1913 -8435
rect 1121 -8549 1154 -8506
rect 1154 -8549 1187 -8506
rect 1088 -8549 1121 -8506
rect 1253 -8549 1286 -8506
rect 1286 -8549 1319 -8506
rect 1220 -8549 1253 -8506
rect 1385 -8549 1418 -8506
rect 1418 -8549 1451 -8506
rect 1352 -8549 1385 -8506
rect 1418 -8549 1451 -8506
rect 1451 -8549 1484 -8506
rect 1484 -8549 1517 -8506
rect 1649 -8549 1682 -8506
rect 1682 -8549 1715 -8506
rect 1616 -8549 1649 -8506
rect 1781 -8549 1814 -8506
rect 1814 -8549 1847 -8506
rect 1748 -8549 1781 -8506
rect 1913 -8549 1946 -8506
rect 1946 -8549 1979 -8506
rect 1880 -8549 1913 -8506
rect 1022 -8620 1055 -8577
rect 1055 -8620 1088 -8577
rect 1088 -8620 1121 -8577
rect 1154 -8620 1187 -8577
rect 1187 -8620 1220 -8577
rect 1220 -8620 1253 -8577
rect 1286 -8620 1319 -8577
rect 1319 -8620 1352 -8577
rect 1352 -8620 1385 -8577
rect 1517 -8620 1550 -8577
rect 1550 -8620 1583 -8577
rect 1484 -8620 1517 -8577
rect 1649 -8620 1682 -8577
rect 1682 -8620 1715 -8577
rect 1616 -8620 1649 -8577
rect 1781 -8620 1814 -8577
rect 1814 -8620 1847 -8577
rect 1748 -8620 1781 -8577
rect 1913 -8620 1946 -8577
rect 1946 -8620 1979 -8577
rect 1880 -8620 1913 -8577
rect 1121 -8691 1154 -8648
rect 1154 -8691 1187 -8648
rect 1088 -8691 1121 -8648
rect 1154 -8691 1187 -8648
rect 1187 -8691 1220 -8648
rect 1220 -8691 1253 -8648
rect 1286 -8691 1319 -8648
rect 1319 -8691 1352 -8648
rect 1352 -8691 1385 -8648
rect 1517 -8691 1550 -8648
rect 1550 -8691 1583 -8648
rect 1484 -8691 1517 -8648
rect 1649 -8691 1682 -8648
rect 1682 -8691 1715 -8648
rect 1616 -8691 1649 -8648
rect 1781 -8691 1814 -8648
rect 1814 -8691 1847 -8648
rect 1748 -8691 1781 -8648
rect 1913 -8691 1946 -8648
rect 1946 -8691 1979 -8648
rect 1880 -8691 1913 -8648
rect 1022 -8762 1055 -8719
rect 1055 -8762 1088 -8719
rect 1088 -8762 1121 -8719
rect 1253 -8762 1286 -8719
rect 1286 -8762 1319 -8719
rect 1220 -8762 1253 -8719
rect 1286 -8762 1319 -8719
rect 1319 -8762 1352 -8719
rect 1352 -8762 1385 -8719
rect 1517 -8762 1550 -8719
rect 1550 -8762 1583 -8719
rect 1484 -8762 1517 -8719
rect 1649 -8762 1682 -8719
rect 1682 -8762 1715 -8719
rect 1616 -8762 1649 -8719
rect 1781 -8762 1814 -8719
rect 1814 -8762 1847 -8719
rect 1748 -8762 1781 -8719
rect 1913 -8762 1946 -8719
rect 1946 -8762 1979 -8719
rect 1880 -8762 1913 -8719
rect 1121 -8833 1154 -8790
rect 1154 -8833 1187 -8790
rect 1088 -8833 1121 -8790
rect 1253 -8833 1286 -8790
rect 1286 -8833 1319 -8790
rect 1220 -8833 1253 -8790
rect 1286 -8833 1319 -8790
rect 1319 -8833 1352 -8790
rect 1352 -8833 1385 -8790
rect 1517 -8833 1550 -8790
rect 1550 -8833 1583 -8790
rect 1484 -8833 1517 -8790
rect 1649 -8833 1682 -8790
rect 1682 -8833 1715 -8790
rect 1616 -8833 1649 -8790
rect 1781 -8833 1814 -8790
rect 1814 -8833 1847 -8790
rect 1748 -8833 1781 -8790
rect 1913 -8833 1946 -8790
rect 1946 -8833 1979 -8790
rect 1880 -8833 1913 -8790
rect 1022 -8904 1055 -8861
rect 1055 -8904 1088 -8861
rect 1088 -8904 1121 -8861
rect 1154 -8904 1187 -8861
rect 1187 -8904 1220 -8861
rect 1220 -8904 1253 -8861
rect 1385 -8904 1418 -8861
rect 1418 -8904 1451 -8861
rect 1352 -8904 1385 -8861
rect 1517 -8904 1550 -8861
rect 1550 -8904 1583 -8861
rect 1484 -8904 1517 -8861
rect 1649 -8904 1682 -8861
rect 1682 -8904 1715 -8861
rect 1616 -8904 1649 -8861
rect 1781 -8904 1814 -8861
rect 1814 -8904 1847 -8861
rect 1748 -8904 1781 -8861
rect 1913 -8904 1946 -8861
rect 1946 -8904 1979 -8861
rect 1880 -8904 1913 -8861
rect 1121 -8975 1154 -8932
rect 1154 -8975 1187 -8932
rect 1088 -8975 1121 -8932
rect 1154 -8975 1187 -8932
rect 1187 -8975 1220 -8932
rect 1220 -8975 1253 -8932
rect 1385 -8975 1418 -8932
rect 1418 -8975 1451 -8932
rect 1352 -8975 1385 -8932
rect 1517 -8975 1550 -8932
rect 1550 -8975 1583 -8932
rect 1484 -8975 1517 -8932
rect 1649 -8975 1682 -8932
rect 1682 -8975 1715 -8932
rect 1616 -8975 1649 -8932
rect 1781 -8975 1814 -8932
rect 1814 -8975 1847 -8932
rect 1748 -8975 1781 -8932
rect 1913 -8975 1946 -8932
rect 1946 -8975 1979 -8932
rect 1880 -8975 1913 -8932
rect 1022 -9046 1055 -9003
rect 1055 -9046 1088 -9003
rect 1088 -9046 1121 -9003
rect 1253 -9046 1286 -9003
rect 1286 -9046 1319 -9003
rect 1220 -9046 1253 -9003
rect 1385 -9046 1418 -9003
rect 1418 -9046 1451 -9003
rect 1352 -9046 1385 -9003
rect 1517 -9046 1550 -9003
rect 1550 -9046 1583 -9003
rect 1484 -9046 1517 -9003
rect 1649 -9046 1682 -9003
rect 1682 -9046 1715 -9003
rect 1616 -9046 1649 -9003
rect 1781 -9046 1814 -9003
rect 1814 -9046 1847 -9003
rect 1748 -9046 1781 -9003
rect 1913 -9046 1946 -9003
rect 1946 -9046 1979 -9003
rect 1880 -9046 1913 -9003
rect 1121 -9117 1154 -9074
rect 1154 -9117 1187 -9074
rect 1088 -9117 1121 -9074
rect 1253 -9117 1286 -9074
rect 1286 -9117 1319 -9074
rect 1220 -9117 1253 -9074
rect 1385 -9117 1418 -9074
rect 1418 -9117 1451 -9074
rect 1352 -9117 1385 -9074
rect 1517 -9117 1550 -9074
rect 1550 -9117 1583 -9074
rect 1484 -9117 1517 -9074
rect 1649 -9117 1682 -9074
rect 1682 -9117 1715 -9074
rect 1616 -9117 1649 -9074
rect 1781 -9117 1814 -9074
rect 1814 -9117 1847 -9074
rect 1748 -9117 1781 -9074
rect 1913 -9117 1946 -9074
rect 1946 -9117 1979 -9074
rect 1880 -9117 1913 -9074
rect 0 192 89 235
rect 132 192 221 235
rect 264 192 353 235
rect 396 192 485 235
rect 528 192 617 235
rect 660 192 749 235
rect 792 192 881 235
rect 1065 192 1154 235
rect 1197 192 1286 235
rect 1329 192 1418 235
rect 1461 192 1550 235
rect 1593 192 1682 235
rect 1725 192 1814 235
rect 1857 192 1946 235
<< pdiffc >>
rect -25 -92 -8 -65
rect 41 -92 58 -65
rect 107 -92 124 -65
rect 173 -92 190 -65
rect 239 -92 256 -65
rect 305 -92 322 -65
rect 371 -92 388 -65
rect 437 -92 454 -65
rect 503 -92 520 -65
rect 569 -92 586 -65
rect 635 -92 652 -65
rect 701 -92 718 -65
rect 767 -92 784 -65
rect 833 -92 850 -65
rect 899 -92 916 -65
rect -25 -163 -8 -136
rect 41 -163 58 -136
rect 107 -163 124 -136
rect 173 -163 190 -136
rect 239 -163 256 -136
rect 305 -163 322 -136
rect 371 -163 388 -136
rect 437 -163 454 -136
rect 503 -163 520 -136
rect 569 -163 586 -136
rect 635 -163 652 -136
rect 701 -163 718 -136
rect 767 -163 784 -136
rect 833 -163 850 -136
rect 899 -163 916 -136
rect -25 -234 -8 -207
rect 41 -234 58 -207
rect 107 -234 124 -207
rect 173 -234 190 -207
rect 239 -234 256 -207
rect 305 -234 322 -207
rect 371 -234 388 -207
rect 437 -234 454 -207
rect 503 -234 520 -207
rect 569 -234 586 -207
rect 635 -234 652 -207
rect 701 -234 718 -207
rect 767 -234 784 -207
rect 833 -234 850 -207
rect 899 -234 916 -207
rect -25 -305 -8 -278
rect 41 -305 58 -278
rect 107 -305 124 -278
rect 173 -305 190 -278
rect 239 -305 256 -278
rect 305 -305 322 -278
rect 371 -305 388 -278
rect 437 -305 454 -278
rect 503 -305 520 -278
rect 569 -305 586 -278
rect 635 -305 652 -278
rect 701 -305 718 -278
rect 767 -305 784 -278
rect 833 -305 850 -278
rect 899 -305 916 -278
rect -25 -376 -8 -349
rect 41 -376 58 -349
rect 107 -376 124 -349
rect 173 -376 190 -349
rect 239 -376 256 -349
rect 305 -376 322 -349
rect 371 -376 388 -349
rect 437 -376 454 -349
rect 503 -376 520 -349
rect 569 -376 586 -349
rect 635 -376 652 -349
rect 701 -376 718 -349
rect 767 -376 784 -349
rect 833 -376 850 -349
rect 899 -376 916 -349
rect -25 -447 -8 -420
rect 41 -447 58 -420
rect 107 -447 124 -420
rect 173 -447 190 -420
rect 239 -447 256 -420
rect 305 -447 322 -420
rect 371 -447 388 -420
rect 437 -447 454 -420
rect 503 -447 520 -420
rect 569 -447 586 -420
rect 635 -447 652 -420
rect 701 -447 718 -420
rect 767 -447 784 -420
rect 833 -447 850 -420
rect 899 -447 916 -420
rect -25 -518 -8 -491
rect 41 -518 58 -491
rect 107 -518 124 -491
rect 173 -518 190 -491
rect 239 -518 256 -491
rect 305 -518 322 -491
rect 371 -518 388 -491
rect 437 -518 454 -491
rect 503 -518 520 -491
rect 569 -518 586 -491
rect 635 -518 652 -491
rect 701 -518 718 -491
rect 767 -518 784 -491
rect 833 -518 850 -491
rect 899 -518 916 -491
rect -25 -589 -8 -562
rect 41 -589 58 -562
rect 107 -589 124 -562
rect 173 -589 190 -562
rect 239 -589 256 -562
rect 305 -589 322 -562
rect 371 -589 388 -562
rect 437 -589 454 -562
rect 503 -589 520 -562
rect 569 -589 586 -562
rect 635 -589 652 -562
rect 701 -589 718 -562
rect 767 -589 784 -562
rect 833 -589 850 -562
rect 899 -589 916 -562
rect -25 -660 -8 -633
rect 41 -660 58 -633
rect 107 -660 124 -633
rect 173 -660 190 -633
rect 239 -660 256 -633
rect 305 -660 322 -633
rect 371 -660 388 -633
rect 437 -660 454 -633
rect 503 -660 520 -633
rect 569 -660 586 -633
rect 635 -660 652 -633
rect 701 -660 718 -633
rect 767 -660 784 -633
rect 833 -660 850 -633
rect 899 -660 916 -633
rect -25 -731 -8 -704
rect 41 -731 58 -704
rect 107 -731 124 -704
rect 173 -731 190 -704
rect 239 -731 256 -704
rect 305 -731 322 -704
rect 371 -731 388 -704
rect 437 -731 454 -704
rect 503 -731 520 -704
rect 569 -731 586 -704
rect 635 -731 652 -704
rect 701 -731 718 -704
rect 767 -731 784 -704
rect 833 -731 850 -704
rect 899 -731 916 -704
rect -25 -802 -8 -775
rect 41 -802 58 -775
rect 107 -802 124 -775
rect 173 -802 190 -775
rect 239 -802 256 -775
rect 305 -802 322 -775
rect 371 -802 388 -775
rect 437 -802 454 -775
rect 503 -802 520 -775
rect 569 -802 586 -775
rect 635 -802 652 -775
rect 701 -802 718 -775
rect 767 -802 784 -775
rect 833 -802 850 -775
rect 899 -802 916 -775
rect -25 -873 -8 -846
rect 41 -873 58 -846
rect 107 -873 124 -846
rect 173 -873 190 -846
rect 239 -873 256 -846
rect 305 -873 322 -846
rect 371 -873 388 -846
rect 437 -873 454 -846
rect 503 -873 520 -846
rect 569 -873 586 -846
rect 635 -873 652 -846
rect 701 -873 718 -846
rect 767 -873 784 -846
rect 833 -873 850 -846
rect 899 -873 916 -846
rect -25 -944 -8 -917
rect 41 -944 58 -917
rect 107 -944 124 -917
rect 173 -944 190 -917
rect 239 -944 256 -917
rect 305 -944 322 -917
rect 371 -944 388 -917
rect 437 -944 454 -917
rect 503 -944 520 -917
rect 569 -944 586 -917
rect 635 -944 652 -917
rect 701 -944 718 -917
rect 767 -944 784 -917
rect 833 -944 850 -917
rect 899 -944 916 -917
rect -25 -1015 -8 -988
rect 41 -1015 58 -988
rect 107 -1015 124 -988
rect 173 -1015 190 -988
rect 239 -1015 256 -988
rect 305 -1015 322 -988
rect 371 -1015 388 -988
rect 437 -1015 454 -988
rect 503 -1015 520 -988
rect 569 -1015 586 -988
rect 635 -1015 652 -988
rect 701 -1015 718 -988
rect 767 -1015 784 -988
rect 833 -1015 850 -988
rect 899 -1015 916 -988
rect -25 -1086 -8 -1059
rect 41 -1086 58 -1059
rect 107 -1086 124 -1059
rect 173 -1086 190 -1059
rect 239 -1086 256 -1059
rect 305 -1086 322 -1059
rect 371 -1086 388 -1059
rect 437 -1086 454 -1059
rect 503 -1086 520 -1059
rect 569 -1086 586 -1059
rect 635 -1086 652 -1059
rect 701 -1086 718 -1059
rect 767 -1086 784 -1059
rect 833 -1086 850 -1059
rect 899 -1086 916 -1059
rect -25 -1157 -8 -1130
rect 41 -1157 58 -1130
rect 107 -1157 124 -1130
rect 173 -1157 190 -1130
rect 239 -1157 256 -1130
rect 305 -1157 322 -1130
rect 371 -1157 388 -1130
rect 437 -1157 454 -1130
rect 503 -1157 520 -1130
rect 569 -1157 586 -1130
rect 635 -1157 652 -1130
rect 701 -1157 718 -1130
rect 767 -1157 784 -1130
rect 833 -1157 850 -1130
rect 899 -1157 916 -1130
rect -25 -1228 -8 -1201
rect 41 -1228 58 -1201
rect 107 -1228 124 -1201
rect 173 -1228 190 -1201
rect 239 -1228 256 -1201
rect 305 -1228 322 -1201
rect 371 -1228 388 -1201
rect 437 -1228 454 -1201
rect 503 -1228 520 -1201
rect 569 -1228 586 -1201
rect 635 -1228 652 -1201
rect 701 -1228 718 -1201
rect 767 -1228 784 -1201
rect 833 -1228 850 -1201
rect 899 -1228 916 -1201
rect -25 -1299 -8 -1272
rect 41 -1299 58 -1272
rect 107 -1299 124 -1272
rect 173 -1299 190 -1272
rect 239 -1299 256 -1272
rect 305 -1299 322 -1272
rect 371 -1299 388 -1272
rect 437 -1299 454 -1272
rect 503 -1299 520 -1272
rect 569 -1299 586 -1272
rect 635 -1299 652 -1272
rect 701 -1299 718 -1272
rect 767 -1299 784 -1272
rect 833 -1299 850 -1272
rect 899 -1299 916 -1272
rect -25 -1370 -8 -1343
rect 41 -1370 58 -1343
rect 107 -1370 124 -1343
rect 173 -1370 190 -1343
rect 239 -1370 256 -1343
rect 305 -1370 322 -1343
rect 371 -1370 388 -1343
rect 437 -1370 454 -1343
rect 503 -1370 520 -1343
rect 569 -1370 586 -1343
rect 635 -1370 652 -1343
rect 701 -1370 718 -1343
rect 767 -1370 784 -1343
rect 833 -1370 850 -1343
rect 899 -1370 916 -1343
rect -25 -1441 -8 -1414
rect 41 -1441 58 -1414
rect 107 -1441 124 -1414
rect 173 -1441 190 -1414
rect 239 -1441 256 -1414
rect 305 -1441 322 -1414
rect 371 -1441 388 -1414
rect 437 -1441 454 -1414
rect 503 -1441 520 -1414
rect 569 -1441 586 -1414
rect 635 -1441 652 -1414
rect 701 -1441 718 -1414
rect 767 -1441 784 -1414
rect 833 -1441 850 -1414
rect 899 -1441 916 -1414
rect -25 -1512 -8 -1485
rect 41 -1512 58 -1485
rect 107 -1512 124 -1485
rect 173 -1512 190 -1485
rect 239 -1512 256 -1485
rect 305 -1512 322 -1485
rect 371 -1512 388 -1485
rect 437 -1512 454 -1485
rect 503 -1512 520 -1485
rect 569 -1512 586 -1485
rect 635 -1512 652 -1485
rect 701 -1512 718 -1485
rect 767 -1512 784 -1485
rect 833 -1512 850 -1485
rect 899 -1512 916 -1485
rect -25 -1583 -8 -1556
rect 41 -1583 58 -1556
rect 107 -1583 124 -1556
rect 173 -1583 190 -1556
rect 239 -1583 256 -1556
rect 305 -1583 322 -1556
rect 371 -1583 388 -1556
rect 437 -1583 454 -1556
rect 503 -1583 520 -1556
rect 569 -1583 586 -1556
rect 635 -1583 652 -1556
rect 701 -1583 718 -1556
rect 767 -1583 784 -1556
rect 833 -1583 850 -1556
rect 899 -1583 916 -1556
rect -25 -1654 -8 -1627
rect 41 -1654 58 -1627
rect 107 -1654 124 -1627
rect 173 -1654 190 -1627
rect 239 -1654 256 -1627
rect 305 -1654 322 -1627
rect 371 -1654 388 -1627
rect 437 -1654 454 -1627
rect 503 -1654 520 -1627
rect 569 -1654 586 -1627
rect 635 -1654 652 -1627
rect 701 -1654 718 -1627
rect 767 -1654 784 -1627
rect 833 -1654 850 -1627
rect 899 -1654 916 -1627
rect -25 -1725 -8 -1698
rect 41 -1725 58 -1698
rect 107 -1725 124 -1698
rect 173 -1725 190 -1698
rect 239 -1725 256 -1698
rect 305 -1725 322 -1698
rect 371 -1725 388 -1698
rect 437 -1725 454 -1698
rect 503 -1725 520 -1698
rect 569 -1725 586 -1698
rect 635 -1725 652 -1698
rect 701 -1725 718 -1698
rect 767 -1725 784 -1698
rect 833 -1725 850 -1698
rect 899 -1725 916 -1698
rect -25 -1796 -8 -1769
rect 41 -1796 58 -1769
rect 107 -1796 124 -1769
rect 173 -1796 190 -1769
rect 239 -1796 256 -1769
rect 305 -1796 322 -1769
rect 371 -1796 388 -1769
rect 437 -1796 454 -1769
rect 503 -1796 520 -1769
rect 569 -1796 586 -1769
rect 635 -1796 652 -1769
rect 701 -1796 718 -1769
rect 767 -1796 784 -1769
rect 833 -1796 850 -1769
rect 899 -1796 916 -1769
rect -25 -1867 -8 -1840
rect 41 -1867 58 -1840
rect 107 -1867 124 -1840
rect 173 -1867 190 -1840
rect 239 -1867 256 -1840
rect 305 -1867 322 -1840
rect 371 -1867 388 -1840
rect 437 -1867 454 -1840
rect 503 -1867 520 -1840
rect 569 -1867 586 -1840
rect 635 -1867 652 -1840
rect 701 -1867 718 -1840
rect 767 -1867 784 -1840
rect 833 -1867 850 -1840
rect 899 -1867 916 -1840
rect -25 -1938 -8 -1911
rect 41 -1938 58 -1911
rect 107 -1938 124 -1911
rect 173 -1938 190 -1911
rect 239 -1938 256 -1911
rect 305 -1938 322 -1911
rect 371 -1938 388 -1911
rect 437 -1938 454 -1911
rect 503 -1938 520 -1911
rect 569 -1938 586 -1911
rect 635 -1938 652 -1911
rect 701 -1938 718 -1911
rect 767 -1938 784 -1911
rect 833 -1938 850 -1911
rect 899 -1938 916 -1911
rect -25 -2009 -8 -1982
rect 41 -2009 58 -1982
rect 107 -2009 124 -1982
rect 173 -2009 190 -1982
rect 239 -2009 256 -1982
rect 305 -2009 322 -1982
rect 371 -2009 388 -1982
rect 437 -2009 454 -1982
rect 503 -2009 520 -1982
rect 569 -2009 586 -1982
rect 635 -2009 652 -1982
rect 701 -2009 718 -1982
rect 767 -2009 784 -1982
rect 833 -2009 850 -1982
rect 899 -2009 916 -1982
rect -25 -2080 -8 -2053
rect 41 -2080 58 -2053
rect 107 -2080 124 -2053
rect 173 -2080 190 -2053
rect 239 -2080 256 -2053
rect 305 -2080 322 -2053
rect 371 -2080 388 -2053
rect 437 -2080 454 -2053
rect 503 -2080 520 -2053
rect 569 -2080 586 -2053
rect 635 -2080 652 -2053
rect 701 -2080 718 -2053
rect 767 -2080 784 -2053
rect 833 -2080 850 -2053
rect 899 -2080 916 -2053
rect -25 -2151 -8 -2124
rect 41 -2151 58 -2124
rect 107 -2151 124 -2124
rect 173 -2151 190 -2124
rect 239 -2151 256 -2124
rect 305 -2151 322 -2124
rect 371 -2151 388 -2124
rect 437 -2151 454 -2124
rect 503 -2151 520 -2124
rect 569 -2151 586 -2124
rect 635 -2151 652 -2124
rect 701 -2151 718 -2124
rect 767 -2151 784 -2124
rect 833 -2151 850 -2124
rect 899 -2151 916 -2124
rect -25 -2222 -8 -2195
rect 41 -2222 58 -2195
rect 107 -2222 124 -2195
rect 173 -2222 190 -2195
rect 239 -2222 256 -2195
rect 305 -2222 322 -2195
rect 371 -2222 388 -2195
rect 437 -2222 454 -2195
rect 503 -2222 520 -2195
rect 569 -2222 586 -2195
rect 635 -2222 652 -2195
rect 701 -2222 718 -2195
rect 767 -2222 784 -2195
rect 833 -2222 850 -2195
rect 899 -2222 916 -2195
rect -25 -2293 -8 -2266
rect 41 -2293 58 -2266
rect 107 -2293 124 -2266
rect 173 -2293 190 -2266
rect 239 -2293 256 -2266
rect 305 -2293 322 -2266
rect 371 -2293 388 -2266
rect 437 -2293 454 -2266
rect 503 -2293 520 -2266
rect 569 -2293 586 -2266
rect 635 -2293 652 -2266
rect 701 -2293 718 -2266
rect 767 -2293 784 -2266
rect 833 -2293 850 -2266
rect 899 -2293 916 -2266
rect -25 -2364 -8 -2337
rect 41 -2364 58 -2337
rect 107 -2364 124 -2337
rect 173 -2364 190 -2337
rect 239 -2364 256 -2337
rect 305 -2364 322 -2337
rect 371 -2364 388 -2337
rect 437 -2364 454 -2337
rect 503 -2364 520 -2337
rect 569 -2364 586 -2337
rect 635 -2364 652 -2337
rect 701 -2364 718 -2337
rect 767 -2364 784 -2337
rect 833 -2364 850 -2337
rect 899 -2364 916 -2337
rect -25 -2435 -8 -2408
rect 41 -2435 58 -2408
rect 107 -2435 124 -2408
rect 173 -2435 190 -2408
rect 239 -2435 256 -2408
rect 305 -2435 322 -2408
rect 371 -2435 388 -2408
rect 437 -2435 454 -2408
rect 503 -2435 520 -2408
rect 569 -2435 586 -2408
rect 635 -2435 652 -2408
rect 701 -2435 718 -2408
rect 767 -2435 784 -2408
rect 833 -2435 850 -2408
rect 899 -2435 916 -2408
rect -25 -2506 -8 -2479
rect 41 -2506 58 -2479
rect 107 -2506 124 -2479
rect 173 -2506 190 -2479
rect 239 -2506 256 -2479
rect 305 -2506 322 -2479
rect 371 -2506 388 -2479
rect 437 -2506 454 -2479
rect 503 -2506 520 -2479
rect 569 -2506 586 -2479
rect 635 -2506 652 -2479
rect 701 -2506 718 -2479
rect 767 -2506 784 -2479
rect 833 -2506 850 -2479
rect 899 -2506 916 -2479
rect -25 -2577 -8 -2550
rect 41 -2577 58 -2550
rect 107 -2577 124 -2550
rect 173 -2577 190 -2550
rect 239 -2577 256 -2550
rect 305 -2577 322 -2550
rect 371 -2577 388 -2550
rect 437 -2577 454 -2550
rect 503 -2577 520 -2550
rect 569 -2577 586 -2550
rect 635 -2577 652 -2550
rect 701 -2577 718 -2550
rect 767 -2577 784 -2550
rect 833 -2577 850 -2550
rect 899 -2577 916 -2550
rect -25 -2648 -8 -2621
rect 41 -2648 58 -2621
rect 107 -2648 124 -2621
rect 173 -2648 190 -2621
rect 239 -2648 256 -2621
rect 305 -2648 322 -2621
rect 371 -2648 388 -2621
rect 437 -2648 454 -2621
rect 503 -2648 520 -2621
rect 569 -2648 586 -2621
rect 635 -2648 652 -2621
rect 701 -2648 718 -2621
rect 767 -2648 784 -2621
rect 833 -2648 850 -2621
rect 899 -2648 916 -2621
rect -25 -2719 -8 -2692
rect 41 -2719 58 -2692
rect 107 -2719 124 -2692
rect 173 -2719 190 -2692
rect 239 -2719 256 -2692
rect 305 -2719 322 -2692
rect 371 -2719 388 -2692
rect 437 -2719 454 -2692
rect 503 -2719 520 -2692
rect 569 -2719 586 -2692
rect 635 -2719 652 -2692
rect 701 -2719 718 -2692
rect 767 -2719 784 -2692
rect 833 -2719 850 -2692
rect 899 -2719 916 -2692
rect -25 -2790 -8 -2763
rect 41 -2790 58 -2763
rect 107 -2790 124 -2763
rect 173 -2790 190 -2763
rect 239 -2790 256 -2763
rect 305 -2790 322 -2763
rect 371 -2790 388 -2763
rect 437 -2790 454 -2763
rect 503 -2790 520 -2763
rect 569 -2790 586 -2763
rect 635 -2790 652 -2763
rect 701 -2790 718 -2763
rect 767 -2790 784 -2763
rect 833 -2790 850 -2763
rect 899 -2790 916 -2763
rect -25 -2861 -8 -2834
rect 41 -2861 58 -2834
rect 107 -2861 124 -2834
rect 173 -2861 190 -2834
rect 239 -2861 256 -2834
rect 305 -2861 322 -2834
rect 371 -2861 388 -2834
rect 437 -2861 454 -2834
rect 503 -2861 520 -2834
rect 569 -2861 586 -2834
rect 635 -2861 652 -2834
rect 701 -2861 718 -2834
rect 767 -2861 784 -2834
rect 833 -2861 850 -2834
rect 899 -2861 916 -2834
rect -25 -2932 -8 -2905
rect 41 -2932 58 -2905
rect 107 -2932 124 -2905
rect 173 -2932 190 -2905
rect 239 -2932 256 -2905
rect 305 -2932 322 -2905
rect 371 -2932 388 -2905
rect 437 -2932 454 -2905
rect 503 -2932 520 -2905
rect 569 -2932 586 -2905
rect 635 -2932 652 -2905
rect 701 -2932 718 -2905
rect 767 -2932 784 -2905
rect 833 -2932 850 -2905
rect 899 -2932 916 -2905
rect -25 -3003 -8 -2976
rect 41 -3003 58 -2976
rect 107 -3003 124 -2976
rect 173 -3003 190 -2976
rect 239 -3003 256 -2976
rect 305 -3003 322 -2976
rect 371 -3003 388 -2976
rect 437 -3003 454 -2976
rect 503 -3003 520 -2976
rect 569 -3003 586 -2976
rect 635 -3003 652 -2976
rect 701 -3003 718 -2976
rect 767 -3003 784 -2976
rect 833 -3003 850 -2976
rect 899 -3003 916 -2976
rect -25 -3074 -8 -3047
rect 41 -3074 58 -3047
rect 107 -3074 124 -3047
rect 173 -3074 190 -3047
rect 239 -3074 256 -3047
rect 305 -3074 322 -3047
rect 371 -3074 388 -3047
rect 437 -3074 454 -3047
rect 503 -3074 520 -3047
rect 569 -3074 586 -3047
rect 635 -3074 652 -3047
rect 701 -3074 718 -3047
rect 767 -3074 784 -3047
rect 833 -3074 850 -3047
rect 899 -3074 916 -3047
rect -25 -3145 -8 -3118
rect 41 -3145 58 -3118
rect 107 -3145 124 -3118
rect 173 -3145 190 -3118
rect 239 -3145 256 -3118
rect 305 -3145 322 -3118
rect 371 -3145 388 -3118
rect 437 -3145 454 -3118
rect 503 -3145 520 -3118
rect 569 -3145 586 -3118
rect 635 -3145 652 -3118
rect 701 -3145 718 -3118
rect 767 -3145 784 -3118
rect 833 -3145 850 -3118
rect 899 -3145 916 -3118
rect -25 -3216 -8 -3189
rect 41 -3216 58 -3189
rect 107 -3216 124 -3189
rect 173 -3216 190 -3189
rect 239 -3216 256 -3189
rect 305 -3216 322 -3189
rect 371 -3216 388 -3189
rect 437 -3216 454 -3189
rect 503 -3216 520 -3189
rect 569 -3216 586 -3189
rect 635 -3216 652 -3189
rect 701 -3216 718 -3189
rect 767 -3216 784 -3189
rect 833 -3216 850 -3189
rect 899 -3216 916 -3189
rect -25 -3287 -8 -3260
rect 41 -3287 58 -3260
rect 107 -3287 124 -3260
rect 173 -3287 190 -3260
rect 239 -3287 256 -3260
rect 305 -3287 322 -3260
rect 371 -3287 388 -3260
rect 437 -3287 454 -3260
rect 503 -3287 520 -3260
rect 569 -3287 586 -3260
rect 635 -3287 652 -3260
rect 701 -3287 718 -3260
rect 767 -3287 784 -3260
rect 833 -3287 850 -3260
rect 899 -3287 916 -3260
rect -25 -3358 -8 -3331
rect 41 -3358 58 -3331
rect 107 -3358 124 -3331
rect 173 -3358 190 -3331
rect 239 -3358 256 -3331
rect 305 -3358 322 -3331
rect 371 -3358 388 -3331
rect 437 -3358 454 -3331
rect 503 -3358 520 -3331
rect 569 -3358 586 -3331
rect 635 -3358 652 -3331
rect 701 -3358 718 -3331
rect 767 -3358 784 -3331
rect 833 -3358 850 -3331
rect 899 -3358 916 -3331
rect -25 -3429 -8 -3402
rect 41 -3429 58 -3402
rect 107 -3429 124 -3402
rect 173 -3429 190 -3402
rect 239 -3429 256 -3402
rect 305 -3429 322 -3402
rect 371 -3429 388 -3402
rect 437 -3429 454 -3402
rect 503 -3429 520 -3402
rect 569 -3429 586 -3402
rect 635 -3429 652 -3402
rect 701 -3429 718 -3402
rect 767 -3429 784 -3402
rect 833 -3429 850 -3402
rect 899 -3429 916 -3402
rect -25 -3500 -8 -3473
rect 41 -3500 58 -3473
rect 107 -3500 124 -3473
rect 173 -3500 190 -3473
rect 239 -3500 256 -3473
rect 305 -3500 322 -3473
rect 371 -3500 388 -3473
rect 437 -3500 454 -3473
rect 503 -3500 520 -3473
rect 569 -3500 586 -3473
rect 635 -3500 652 -3473
rect 701 -3500 718 -3473
rect 767 -3500 784 -3473
rect 833 -3500 850 -3473
rect 899 -3500 916 -3473
rect -25 -3571 -8 -3544
rect 41 -3571 58 -3544
rect 107 -3571 124 -3544
rect 173 -3571 190 -3544
rect 239 -3571 256 -3544
rect 305 -3571 322 -3544
rect 371 -3571 388 -3544
rect 437 -3571 454 -3544
rect 503 -3571 520 -3544
rect 569 -3571 586 -3544
rect 635 -3571 652 -3544
rect 701 -3571 718 -3544
rect 767 -3571 784 -3544
rect 833 -3571 850 -3544
rect 899 -3571 916 -3544
rect -25 -3642 -8 -3615
rect 41 -3642 58 -3615
rect 107 -3642 124 -3615
rect 173 -3642 190 -3615
rect 239 -3642 256 -3615
rect 305 -3642 322 -3615
rect 371 -3642 388 -3615
rect 437 -3642 454 -3615
rect 503 -3642 520 -3615
rect 569 -3642 586 -3615
rect 635 -3642 652 -3615
rect 701 -3642 718 -3615
rect 767 -3642 784 -3615
rect 833 -3642 850 -3615
rect 899 -3642 916 -3615
rect -25 -3713 -8 -3686
rect 41 -3713 58 -3686
rect 107 -3713 124 -3686
rect 173 -3713 190 -3686
rect 239 -3713 256 -3686
rect 305 -3713 322 -3686
rect 371 -3713 388 -3686
rect 437 -3713 454 -3686
rect 503 -3713 520 -3686
rect 569 -3713 586 -3686
rect 635 -3713 652 -3686
rect 701 -3713 718 -3686
rect 767 -3713 784 -3686
rect 833 -3713 850 -3686
rect 899 -3713 916 -3686
rect -25 -3784 -8 -3757
rect 41 -3784 58 -3757
rect 107 -3784 124 -3757
rect 173 -3784 190 -3757
rect 239 -3784 256 -3757
rect 305 -3784 322 -3757
rect 371 -3784 388 -3757
rect 437 -3784 454 -3757
rect 503 -3784 520 -3757
rect 569 -3784 586 -3757
rect 635 -3784 652 -3757
rect 701 -3784 718 -3757
rect 767 -3784 784 -3757
rect 833 -3784 850 -3757
rect 899 -3784 916 -3757
rect -25 -3855 -8 -3828
rect 41 -3855 58 -3828
rect 107 -3855 124 -3828
rect 173 -3855 190 -3828
rect 239 -3855 256 -3828
rect 305 -3855 322 -3828
rect 371 -3855 388 -3828
rect 437 -3855 454 -3828
rect 503 -3855 520 -3828
rect 569 -3855 586 -3828
rect 635 -3855 652 -3828
rect 701 -3855 718 -3828
rect 767 -3855 784 -3828
rect 833 -3855 850 -3828
rect 899 -3855 916 -3828
rect -25 -3926 -8 -3899
rect 41 -3926 58 -3899
rect 107 -3926 124 -3899
rect 173 -3926 190 -3899
rect 239 -3926 256 -3899
rect 305 -3926 322 -3899
rect 371 -3926 388 -3899
rect 437 -3926 454 -3899
rect 503 -3926 520 -3899
rect 569 -3926 586 -3899
rect 635 -3926 652 -3899
rect 701 -3926 718 -3899
rect 767 -3926 784 -3899
rect 833 -3926 850 -3899
rect 899 -3926 916 -3899
rect -25 -3997 -8 -3970
rect 41 -3997 58 -3970
rect 107 -3997 124 -3970
rect 173 -3997 190 -3970
rect 239 -3997 256 -3970
rect 305 -3997 322 -3970
rect 371 -3997 388 -3970
rect 437 -3997 454 -3970
rect 503 -3997 520 -3970
rect 569 -3997 586 -3970
rect 635 -3997 652 -3970
rect 701 -3997 718 -3970
rect 767 -3997 784 -3970
rect 833 -3997 850 -3970
rect 899 -3997 916 -3970
rect -25 -4068 -8 -4041
rect 41 -4068 58 -4041
rect 107 -4068 124 -4041
rect 173 -4068 190 -4041
rect 239 -4068 256 -4041
rect 305 -4068 322 -4041
rect 371 -4068 388 -4041
rect 437 -4068 454 -4041
rect 503 -4068 520 -4041
rect 569 -4068 586 -4041
rect 635 -4068 652 -4041
rect 701 -4068 718 -4041
rect 767 -4068 784 -4041
rect 833 -4068 850 -4041
rect 899 -4068 916 -4041
rect -25 -4139 -8 -4112
rect 41 -4139 58 -4112
rect 107 -4139 124 -4112
rect 173 -4139 190 -4112
rect 239 -4139 256 -4112
rect 305 -4139 322 -4112
rect 371 -4139 388 -4112
rect 437 -4139 454 -4112
rect 503 -4139 520 -4112
rect 569 -4139 586 -4112
rect 635 -4139 652 -4112
rect 701 -4139 718 -4112
rect 767 -4139 784 -4112
rect 833 -4139 850 -4112
rect 899 -4139 916 -4112
rect -25 -4210 -8 -4183
rect 41 -4210 58 -4183
rect 107 -4210 124 -4183
rect 173 -4210 190 -4183
rect 239 -4210 256 -4183
rect 305 -4210 322 -4183
rect 371 -4210 388 -4183
rect 437 -4210 454 -4183
rect 503 -4210 520 -4183
rect 569 -4210 586 -4183
rect 635 -4210 652 -4183
rect 701 -4210 718 -4183
rect 767 -4210 784 -4183
rect 833 -4210 850 -4183
rect 899 -4210 916 -4183
rect -25 -4281 -8 -4254
rect 41 -4281 58 -4254
rect 107 -4281 124 -4254
rect 173 -4281 190 -4254
rect 239 -4281 256 -4254
rect 305 -4281 322 -4254
rect 371 -4281 388 -4254
rect 437 -4281 454 -4254
rect 503 -4281 520 -4254
rect 569 -4281 586 -4254
rect 635 -4281 652 -4254
rect 701 -4281 718 -4254
rect 767 -4281 784 -4254
rect 833 -4281 850 -4254
rect 899 -4281 916 -4254
rect -25 -4352 -8 -4325
rect 41 -4352 58 -4325
rect 107 -4352 124 -4325
rect 173 -4352 190 -4325
rect 239 -4352 256 -4325
rect 305 -4352 322 -4325
rect 371 -4352 388 -4325
rect 437 -4352 454 -4325
rect 503 -4352 520 -4325
rect 569 -4352 586 -4325
rect 635 -4352 652 -4325
rect 701 -4352 718 -4325
rect 767 -4352 784 -4325
rect 833 -4352 850 -4325
rect 899 -4352 916 -4325
rect -25 -4423 -8 -4396
rect 41 -4423 58 -4396
rect 107 -4423 124 -4396
rect 173 -4423 190 -4396
rect 239 -4423 256 -4396
rect 305 -4423 322 -4396
rect 371 -4423 388 -4396
rect 437 -4423 454 -4396
rect 503 -4423 520 -4396
rect 569 -4423 586 -4396
rect 635 -4423 652 -4396
rect 701 -4423 718 -4396
rect 767 -4423 784 -4396
rect 833 -4423 850 -4396
rect 899 -4423 916 -4396
rect -25 -4494 -8 -4467
rect 41 -4494 58 -4467
rect 107 -4494 124 -4467
rect 173 -4494 190 -4467
rect 239 -4494 256 -4467
rect 305 -4494 322 -4467
rect 371 -4494 388 -4467
rect 437 -4494 454 -4467
rect 503 -4494 520 -4467
rect 569 -4494 586 -4467
rect 635 -4494 652 -4467
rect 701 -4494 718 -4467
rect 767 -4494 784 -4467
rect 833 -4494 850 -4467
rect 899 -4494 916 -4467
rect -25 -4565 -8 -4538
rect 41 -4565 58 -4538
rect 107 -4565 124 -4538
rect 173 -4565 190 -4538
rect 239 -4565 256 -4538
rect 305 -4565 322 -4538
rect 371 -4565 388 -4538
rect 437 -4565 454 -4538
rect 503 -4565 520 -4538
rect 569 -4565 586 -4538
rect 635 -4565 652 -4538
rect 701 -4565 718 -4538
rect 767 -4565 784 -4538
rect 833 -4565 850 -4538
rect 899 -4565 916 -4538
rect -25 -4636 -8 -4609
rect 41 -4636 58 -4609
rect 107 -4636 124 -4609
rect 173 -4636 190 -4609
rect 239 -4636 256 -4609
rect 305 -4636 322 -4609
rect 371 -4636 388 -4609
rect 437 -4636 454 -4609
rect 503 -4636 520 -4609
rect 569 -4636 586 -4609
rect 635 -4636 652 -4609
rect 701 -4636 718 -4609
rect 767 -4636 784 -4609
rect 833 -4636 850 -4609
rect 899 -4636 916 -4609
rect -25 -4707 -8 -4680
rect 41 -4707 58 -4680
rect 107 -4707 124 -4680
rect 173 -4707 190 -4680
rect 239 -4707 256 -4680
rect 305 -4707 322 -4680
rect 371 -4707 388 -4680
rect 437 -4707 454 -4680
rect 503 -4707 520 -4680
rect 569 -4707 586 -4680
rect 635 -4707 652 -4680
rect 701 -4707 718 -4680
rect 767 -4707 784 -4680
rect 833 -4707 850 -4680
rect 899 -4707 916 -4680
rect -25 -4778 -8 -4751
rect 41 -4778 58 -4751
rect 107 -4778 124 -4751
rect 173 -4778 190 -4751
rect 239 -4778 256 -4751
rect 305 -4778 322 -4751
rect 371 -4778 388 -4751
rect 437 -4778 454 -4751
rect 503 -4778 520 -4751
rect 569 -4778 586 -4751
rect 635 -4778 652 -4751
rect 701 -4778 718 -4751
rect 767 -4778 784 -4751
rect 833 -4778 850 -4751
rect 899 -4778 916 -4751
rect -25 -4849 -8 -4822
rect 41 -4849 58 -4822
rect 107 -4849 124 -4822
rect 173 -4849 190 -4822
rect 239 -4849 256 -4822
rect 305 -4849 322 -4822
rect 371 -4849 388 -4822
rect 437 -4849 454 -4822
rect 503 -4849 520 -4822
rect 569 -4849 586 -4822
rect 635 -4849 652 -4822
rect 701 -4849 718 -4822
rect 767 -4849 784 -4822
rect 833 -4849 850 -4822
rect 899 -4849 916 -4822
rect -25 -4920 -8 -4893
rect 41 -4920 58 -4893
rect 107 -4920 124 -4893
rect 173 -4920 190 -4893
rect 239 -4920 256 -4893
rect 305 -4920 322 -4893
rect 371 -4920 388 -4893
rect 437 -4920 454 -4893
rect 503 -4920 520 -4893
rect 569 -4920 586 -4893
rect 635 -4920 652 -4893
rect 701 -4920 718 -4893
rect 767 -4920 784 -4893
rect 833 -4920 850 -4893
rect 899 -4920 916 -4893
rect -25 -4991 -8 -4964
rect 41 -4991 58 -4964
rect 107 -4991 124 -4964
rect 173 -4991 190 -4964
rect 239 -4991 256 -4964
rect 305 -4991 322 -4964
rect 371 -4991 388 -4964
rect 437 -4991 454 -4964
rect 503 -4991 520 -4964
rect 569 -4991 586 -4964
rect 635 -4991 652 -4964
rect 701 -4991 718 -4964
rect 767 -4991 784 -4964
rect 833 -4991 850 -4964
rect 899 -4991 916 -4964
rect -25 -5062 -8 -5035
rect 41 -5062 58 -5035
rect 107 -5062 124 -5035
rect 173 -5062 190 -5035
rect 239 -5062 256 -5035
rect 305 -5062 322 -5035
rect 371 -5062 388 -5035
rect 437 -5062 454 -5035
rect 503 -5062 520 -5035
rect 569 -5062 586 -5035
rect 635 -5062 652 -5035
rect 701 -5062 718 -5035
rect 767 -5062 784 -5035
rect 833 -5062 850 -5035
rect 899 -5062 916 -5035
rect -25 -5133 -8 -5106
rect 41 -5133 58 -5106
rect 107 -5133 124 -5106
rect 173 -5133 190 -5106
rect 239 -5133 256 -5106
rect 305 -5133 322 -5106
rect 371 -5133 388 -5106
rect 437 -5133 454 -5106
rect 503 -5133 520 -5106
rect 569 -5133 586 -5106
rect 635 -5133 652 -5106
rect 701 -5133 718 -5106
rect 767 -5133 784 -5106
rect 833 -5133 850 -5106
rect 899 -5133 916 -5106
rect -25 -5204 -8 -5177
rect 41 -5204 58 -5177
rect 107 -5204 124 -5177
rect 173 -5204 190 -5177
rect 239 -5204 256 -5177
rect 305 -5204 322 -5177
rect 371 -5204 388 -5177
rect 437 -5204 454 -5177
rect 503 -5204 520 -5177
rect 569 -5204 586 -5177
rect 635 -5204 652 -5177
rect 701 -5204 718 -5177
rect 767 -5204 784 -5177
rect 833 -5204 850 -5177
rect 899 -5204 916 -5177
rect -25 -5275 -8 -5248
rect 41 -5275 58 -5248
rect 107 -5275 124 -5248
rect 173 -5275 190 -5248
rect 239 -5275 256 -5248
rect 305 -5275 322 -5248
rect 371 -5275 388 -5248
rect 437 -5275 454 -5248
rect 503 -5275 520 -5248
rect 569 -5275 586 -5248
rect 635 -5275 652 -5248
rect 701 -5275 718 -5248
rect 767 -5275 784 -5248
rect 833 -5275 850 -5248
rect 899 -5275 916 -5248
rect -25 -5346 -8 -5319
rect 41 -5346 58 -5319
rect 107 -5346 124 -5319
rect 173 -5346 190 -5319
rect 239 -5346 256 -5319
rect 305 -5346 322 -5319
rect 371 -5346 388 -5319
rect 437 -5346 454 -5319
rect 503 -5346 520 -5319
rect 569 -5346 586 -5319
rect 635 -5346 652 -5319
rect 701 -5346 718 -5319
rect 767 -5346 784 -5319
rect 833 -5346 850 -5319
rect 899 -5346 916 -5319
rect -25 -5417 -8 -5390
rect 41 -5417 58 -5390
rect 107 -5417 124 -5390
rect 173 -5417 190 -5390
rect 239 -5417 256 -5390
rect 305 -5417 322 -5390
rect 371 -5417 388 -5390
rect 437 -5417 454 -5390
rect 503 -5417 520 -5390
rect 569 -5417 586 -5390
rect 635 -5417 652 -5390
rect 701 -5417 718 -5390
rect 767 -5417 784 -5390
rect 833 -5417 850 -5390
rect 899 -5417 916 -5390
rect -25 -5488 -8 -5461
rect 41 -5488 58 -5461
rect 107 -5488 124 -5461
rect 173 -5488 190 -5461
rect 239 -5488 256 -5461
rect 305 -5488 322 -5461
rect 371 -5488 388 -5461
rect 437 -5488 454 -5461
rect 503 -5488 520 -5461
rect 569 -5488 586 -5461
rect 635 -5488 652 -5461
rect 701 -5488 718 -5461
rect 767 -5488 784 -5461
rect 833 -5488 850 -5461
rect 899 -5488 916 -5461
rect -25 -5559 -8 -5532
rect 41 -5559 58 -5532
rect 107 -5559 124 -5532
rect 173 -5559 190 -5532
rect 239 -5559 256 -5532
rect 305 -5559 322 -5532
rect 371 -5559 388 -5532
rect 437 -5559 454 -5532
rect 503 -5559 520 -5532
rect 569 -5559 586 -5532
rect 635 -5559 652 -5532
rect 701 -5559 718 -5532
rect 767 -5559 784 -5532
rect 833 -5559 850 -5532
rect 899 -5559 916 -5532
rect -25 -5630 -8 -5603
rect 41 -5630 58 -5603
rect 107 -5630 124 -5603
rect 173 -5630 190 -5603
rect 239 -5630 256 -5603
rect 305 -5630 322 -5603
rect 371 -5630 388 -5603
rect 437 -5630 454 -5603
rect 503 -5630 520 -5603
rect 569 -5630 586 -5603
rect 635 -5630 652 -5603
rect 701 -5630 718 -5603
rect 767 -5630 784 -5603
rect 833 -5630 850 -5603
rect 899 -5630 916 -5603
rect -25 -5701 -8 -5674
rect 41 -5701 58 -5674
rect 107 -5701 124 -5674
rect 173 -5701 190 -5674
rect 239 -5701 256 -5674
rect 305 -5701 322 -5674
rect 371 -5701 388 -5674
rect 437 -5701 454 -5674
rect 503 -5701 520 -5674
rect 569 -5701 586 -5674
rect 635 -5701 652 -5674
rect 701 -5701 718 -5674
rect 767 -5701 784 -5674
rect 833 -5701 850 -5674
rect 899 -5701 916 -5674
rect -25 -5772 -8 -5745
rect 41 -5772 58 -5745
rect 107 -5772 124 -5745
rect 173 -5772 190 -5745
rect 239 -5772 256 -5745
rect 305 -5772 322 -5745
rect 371 -5772 388 -5745
rect 437 -5772 454 -5745
rect 503 -5772 520 -5745
rect 569 -5772 586 -5745
rect 635 -5772 652 -5745
rect 701 -5772 718 -5745
rect 767 -5772 784 -5745
rect 833 -5772 850 -5745
rect 899 -5772 916 -5745
rect -25 -5843 -8 -5816
rect 41 -5843 58 -5816
rect 107 -5843 124 -5816
rect 173 -5843 190 -5816
rect 239 -5843 256 -5816
rect 305 -5843 322 -5816
rect 371 -5843 388 -5816
rect 437 -5843 454 -5816
rect 503 -5843 520 -5816
rect 569 -5843 586 -5816
rect 635 -5843 652 -5816
rect 701 -5843 718 -5816
rect 767 -5843 784 -5816
rect 833 -5843 850 -5816
rect 899 -5843 916 -5816
rect -25 -5914 -8 -5887
rect 41 -5914 58 -5887
rect 107 -5914 124 -5887
rect 173 -5914 190 -5887
rect 239 -5914 256 -5887
rect 305 -5914 322 -5887
rect 371 -5914 388 -5887
rect 437 -5914 454 -5887
rect 503 -5914 520 -5887
rect 569 -5914 586 -5887
rect 635 -5914 652 -5887
rect 701 -5914 718 -5887
rect 767 -5914 784 -5887
rect 833 -5914 850 -5887
rect 899 -5914 916 -5887
rect -25 -5985 -8 -5958
rect 41 -5985 58 -5958
rect 107 -5985 124 -5958
rect 173 -5985 190 -5958
rect 239 -5985 256 -5958
rect 305 -5985 322 -5958
rect 371 -5985 388 -5958
rect 437 -5985 454 -5958
rect 503 -5985 520 -5958
rect 569 -5985 586 -5958
rect 635 -5985 652 -5958
rect 701 -5985 718 -5958
rect 767 -5985 784 -5958
rect 833 -5985 850 -5958
rect 899 -5985 916 -5958
rect -25 -6056 -8 -6029
rect 41 -6056 58 -6029
rect 107 -6056 124 -6029
rect 173 -6056 190 -6029
rect 239 -6056 256 -6029
rect 305 -6056 322 -6029
rect 371 -6056 388 -6029
rect 437 -6056 454 -6029
rect 503 -6056 520 -6029
rect 569 -6056 586 -6029
rect 635 -6056 652 -6029
rect 701 -6056 718 -6029
rect 767 -6056 784 -6029
rect 833 -6056 850 -6029
rect 899 -6056 916 -6029
rect -25 -6127 -8 -6100
rect 41 -6127 58 -6100
rect 107 -6127 124 -6100
rect 173 -6127 190 -6100
rect 239 -6127 256 -6100
rect 305 -6127 322 -6100
rect 371 -6127 388 -6100
rect 437 -6127 454 -6100
rect 503 -6127 520 -6100
rect 569 -6127 586 -6100
rect 635 -6127 652 -6100
rect 701 -6127 718 -6100
rect 767 -6127 784 -6100
rect 833 -6127 850 -6100
rect 899 -6127 916 -6100
rect -25 -6198 -8 -6171
rect 41 -6198 58 -6171
rect 107 -6198 124 -6171
rect 173 -6198 190 -6171
rect 239 -6198 256 -6171
rect 305 -6198 322 -6171
rect 371 -6198 388 -6171
rect 437 -6198 454 -6171
rect 503 -6198 520 -6171
rect 569 -6198 586 -6171
rect 635 -6198 652 -6171
rect 701 -6198 718 -6171
rect 767 -6198 784 -6171
rect 833 -6198 850 -6171
rect 899 -6198 916 -6171
rect -25 -6269 -8 -6242
rect 41 -6269 58 -6242
rect 107 -6269 124 -6242
rect 173 -6269 190 -6242
rect 239 -6269 256 -6242
rect 305 -6269 322 -6242
rect 371 -6269 388 -6242
rect 437 -6269 454 -6242
rect 503 -6269 520 -6242
rect 569 -6269 586 -6242
rect 635 -6269 652 -6242
rect 701 -6269 718 -6242
rect 767 -6269 784 -6242
rect 833 -6269 850 -6242
rect 899 -6269 916 -6242
rect -25 -6340 -8 -6313
rect 41 -6340 58 -6313
rect 107 -6340 124 -6313
rect 173 -6340 190 -6313
rect 239 -6340 256 -6313
rect 305 -6340 322 -6313
rect 371 -6340 388 -6313
rect 437 -6340 454 -6313
rect 503 -6340 520 -6313
rect 569 -6340 586 -6313
rect 635 -6340 652 -6313
rect 701 -6340 718 -6313
rect 767 -6340 784 -6313
rect 833 -6340 850 -6313
rect 899 -6340 916 -6313
rect -25 -6411 -8 -6384
rect 41 -6411 58 -6384
rect 107 -6411 124 -6384
rect 173 -6411 190 -6384
rect 239 -6411 256 -6384
rect 305 -6411 322 -6384
rect 371 -6411 388 -6384
rect 437 -6411 454 -6384
rect 503 -6411 520 -6384
rect 569 -6411 586 -6384
rect 635 -6411 652 -6384
rect 701 -6411 718 -6384
rect 767 -6411 784 -6384
rect 833 -6411 850 -6384
rect 899 -6411 916 -6384
rect -25 -6482 -8 -6455
rect 41 -6482 58 -6455
rect 107 -6482 124 -6455
rect 173 -6482 190 -6455
rect 239 -6482 256 -6455
rect 305 -6482 322 -6455
rect 371 -6482 388 -6455
rect 437 -6482 454 -6455
rect 503 -6482 520 -6455
rect 569 -6482 586 -6455
rect 635 -6482 652 -6455
rect 701 -6482 718 -6455
rect 767 -6482 784 -6455
rect 833 -6482 850 -6455
rect 899 -6482 916 -6455
rect -25 -6553 -8 -6526
rect 41 -6553 58 -6526
rect 107 -6553 124 -6526
rect 173 -6553 190 -6526
rect 239 -6553 256 -6526
rect 305 -6553 322 -6526
rect 371 -6553 388 -6526
rect 437 -6553 454 -6526
rect 503 -6553 520 -6526
rect 569 -6553 586 -6526
rect 635 -6553 652 -6526
rect 701 -6553 718 -6526
rect 767 -6553 784 -6526
rect 833 -6553 850 -6526
rect 899 -6553 916 -6526
rect -25 -6624 -8 -6597
rect 41 -6624 58 -6597
rect 107 -6624 124 -6597
rect 173 -6624 190 -6597
rect 239 -6624 256 -6597
rect 305 -6624 322 -6597
rect 371 -6624 388 -6597
rect 437 -6624 454 -6597
rect 503 -6624 520 -6597
rect 569 -6624 586 -6597
rect 635 -6624 652 -6597
rect 701 -6624 718 -6597
rect 767 -6624 784 -6597
rect 833 -6624 850 -6597
rect 899 -6624 916 -6597
rect -25 -6695 -8 -6668
rect 41 -6695 58 -6668
rect 107 -6695 124 -6668
rect 173 -6695 190 -6668
rect 239 -6695 256 -6668
rect 305 -6695 322 -6668
rect 371 -6695 388 -6668
rect 437 -6695 454 -6668
rect 503 -6695 520 -6668
rect 569 -6695 586 -6668
rect 635 -6695 652 -6668
rect 701 -6695 718 -6668
rect 767 -6695 784 -6668
rect 833 -6695 850 -6668
rect 899 -6695 916 -6668
rect -25 -6766 -8 -6739
rect 41 -6766 58 -6739
rect 107 -6766 124 -6739
rect 173 -6766 190 -6739
rect 239 -6766 256 -6739
rect 305 -6766 322 -6739
rect 371 -6766 388 -6739
rect 437 -6766 454 -6739
rect 503 -6766 520 -6739
rect 569 -6766 586 -6739
rect 635 -6766 652 -6739
rect 701 -6766 718 -6739
rect 767 -6766 784 -6739
rect 833 -6766 850 -6739
rect 899 -6766 916 -6739
rect -25 -6837 -8 -6810
rect 41 -6837 58 -6810
rect 107 -6837 124 -6810
rect 173 -6837 190 -6810
rect 239 -6837 256 -6810
rect 305 -6837 322 -6810
rect 371 -6837 388 -6810
rect 437 -6837 454 -6810
rect 503 -6837 520 -6810
rect 569 -6837 586 -6810
rect 635 -6837 652 -6810
rect 701 -6837 718 -6810
rect 767 -6837 784 -6810
rect 833 -6837 850 -6810
rect 899 -6837 916 -6810
rect -25 -6908 -8 -6881
rect 41 -6908 58 -6881
rect 107 -6908 124 -6881
rect 173 -6908 190 -6881
rect 239 -6908 256 -6881
rect 305 -6908 322 -6881
rect 371 -6908 388 -6881
rect 437 -6908 454 -6881
rect 503 -6908 520 -6881
rect 569 -6908 586 -6881
rect 635 -6908 652 -6881
rect 701 -6908 718 -6881
rect 767 -6908 784 -6881
rect 833 -6908 850 -6881
rect 899 -6908 916 -6881
rect -25 -6979 -8 -6952
rect 41 -6979 58 -6952
rect 107 -6979 124 -6952
rect 173 -6979 190 -6952
rect 239 -6979 256 -6952
rect 305 -6979 322 -6952
rect 371 -6979 388 -6952
rect 437 -6979 454 -6952
rect 503 -6979 520 -6952
rect 569 -6979 586 -6952
rect 635 -6979 652 -6952
rect 701 -6979 718 -6952
rect 767 -6979 784 -6952
rect 833 -6979 850 -6952
rect 899 -6979 916 -6952
rect -25 -7050 -8 -7023
rect 41 -7050 58 -7023
rect 107 -7050 124 -7023
rect 173 -7050 190 -7023
rect 239 -7050 256 -7023
rect 305 -7050 322 -7023
rect 371 -7050 388 -7023
rect 437 -7050 454 -7023
rect 503 -7050 520 -7023
rect 569 -7050 586 -7023
rect 635 -7050 652 -7023
rect 701 -7050 718 -7023
rect 767 -7050 784 -7023
rect 833 -7050 850 -7023
rect 899 -7050 916 -7023
rect -25 -7121 -8 -7094
rect 41 -7121 58 -7094
rect 107 -7121 124 -7094
rect 173 -7121 190 -7094
rect 239 -7121 256 -7094
rect 305 -7121 322 -7094
rect 371 -7121 388 -7094
rect 437 -7121 454 -7094
rect 503 -7121 520 -7094
rect 569 -7121 586 -7094
rect 635 -7121 652 -7094
rect 701 -7121 718 -7094
rect 767 -7121 784 -7094
rect 833 -7121 850 -7094
rect 899 -7121 916 -7094
rect -25 -7192 -8 -7165
rect 41 -7192 58 -7165
rect 107 -7192 124 -7165
rect 173 -7192 190 -7165
rect 239 -7192 256 -7165
rect 305 -7192 322 -7165
rect 371 -7192 388 -7165
rect 437 -7192 454 -7165
rect 503 -7192 520 -7165
rect 569 -7192 586 -7165
rect 635 -7192 652 -7165
rect 701 -7192 718 -7165
rect 767 -7192 784 -7165
rect 833 -7192 850 -7165
rect 899 -7192 916 -7165
rect -25 -7263 -8 -7236
rect 41 -7263 58 -7236
rect 107 -7263 124 -7236
rect 173 -7263 190 -7236
rect 239 -7263 256 -7236
rect 305 -7263 322 -7236
rect 371 -7263 388 -7236
rect 437 -7263 454 -7236
rect 503 -7263 520 -7236
rect 569 -7263 586 -7236
rect 635 -7263 652 -7236
rect 701 -7263 718 -7236
rect 767 -7263 784 -7236
rect 833 -7263 850 -7236
rect 899 -7263 916 -7236
rect -25 -7334 -8 -7307
rect 41 -7334 58 -7307
rect 107 -7334 124 -7307
rect 173 -7334 190 -7307
rect 239 -7334 256 -7307
rect 305 -7334 322 -7307
rect 371 -7334 388 -7307
rect 437 -7334 454 -7307
rect 503 -7334 520 -7307
rect 569 -7334 586 -7307
rect 635 -7334 652 -7307
rect 701 -7334 718 -7307
rect 767 -7334 784 -7307
rect 833 -7334 850 -7307
rect 899 -7334 916 -7307
rect -25 -7405 -8 -7378
rect 41 -7405 58 -7378
rect 107 -7405 124 -7378
rect 173 -7405 190 -7378
rect 239 -7405 256 -7378
rect 305 -7405 322 -7378
rect 371 -7405 388 -7378
rect 437 -7405 454 -7378
rect 503 -7405 520 -7378
rect 569 -7405 586 -7378
rect 635 -7405 652 -7378
rect 701 -7405 718 -7378
rect 767 -7405 784 -7378
rect 833 -7405 850 -7378
rect 899 -7405 916 -7378
rect -25 -7476 -8 -7449
rect 41 -7476 58 -7449
rect 107 -7476 124 -7449
rect 173 -7476 190 -7449
rect 239 -7476 256 -7449
rect 305 -7476 322 -7449
rect 371 -7476 388 -7449
rect 437 -7476 454 -7449
rect 503 -7476 520 -7449
rect 569 -7476 586 -7449
rect 635 -7476 652 -7449
rect 701 -7476 718 -7449
rect 767 -7476 784 -7449
rect 833 -7476 850 -7449
rect 899 -7476 916 -7449
rect -25 -7547 -8 -7520
rect 41 -7547 58 -7520
rect 107 -7547 124 -7520
rect 173 -7547 190 -7520
rect 239 -7547 256 -7520
rect 305 -7547 322 -7520
rect 371 -7547 388 -7520
rect 437 -7547 454 -7520
rect 503 -7547 520 -7520
rect 569 -7547 586 -7520
rect 635 -7547 652 -7520
rect 701 -7547 718 -7520
rect 767 -7547 784 -7520
rect 833 -7547 850 -7520
rect 899 -7547 916 -7520
rect -25 -7618 -8 -7591
rect 41 -7618 58 -7591
rect 107 -7618 124 -7591
rect 173 -7618 190 -7591
rect 239 -7618 256 -7591
rect 305 -7618 322 -7591
rect 371 -7618 388 -7591
rect 437 -7618 454 -7591
rect 503 -7618 520 -7591
rect 569 -7618 586 -7591
rect 635 -7618 652 -7591
rect 701 -7618 718 -7591
rect 767 -7618 784 -7591
rect 833 -7618 850 -7591
rect 899 -7618 916 -7591
rect -25 -7689 -8 -7662
rect 41 -7689 58 -7662
rect 107 -7689 124 -7662
rect 173 -7689 190 -7662
rect 239 -7689 256 -7662
rect 305 -7689 322 -7662
rect 371 -7689 388 -7662
rect 437 -7689 454 -7662
rect 503 -7689 520 -7662
rect 569 -7689 586 -7662
rect 635 -7689 652 -7662
rect 701 -7689 718 -7662
rect 767 -7689 784 -7662
rect 833 -7689 850 -7662
rect 899 -7689 916 -7662
rect -25 -7760 -8 -7733
rect 41 -7760 58 -7733
rect 107 -7760 124 -7733
rect 173 -7760 190 -7733
rect 239 -7760 256 -7733
rect 305 -7760 322 -7733
rect 371 -7760 388 -7733
rect 437 -7760 454 -7733
rect 503 -7760 520 -7733
rect 569 -7760 586 -7733
rect 635 -7760 652 -7733
rect 701 -7760 718 -7733
rect 767 -7760 784 -7733
rect 833 -7760 850 -7733
rect 899 -7760 916 -7733
rect -25 -7831 -8 -7804
rect 41 -7831 58 -7804
rect 107 -7831 124 -7804
rect 173 -7831 190 -7804
rect 239 -7831 256 -7804
rect 305 -7831 322 -7804
rect 371 -7831 388 -7804
rect 437 -7831 454 -7804
rect 503 -7831 520 -7804
rect 569 -7831 586 -7804
rect 635 -7831 652 -7804
rect 701 -7831 718 -7804
rect 767 -7831 784 -7804
rect 833 -7831 850 -7804
rect 899 -7831 916 -7804
rect -25 -7902 -8 -7875
rect 41 -7902 58 -7875
rect 107 -7902 124 -7875
rect 173 -7902 190 -7875
rect 239 -7902 256 -7875
rect 305 -7902 322 -7875
rect 371 -7902 388 -7875
rect 437 -7902 454 -7875
rect 503 -7902 520 -7875
rect 569 -7902 586 -7875
rect 635 -7902 652 -7875
rect 701 -7902 718 -7875
rect 767 -7902 784 -7875
rect 833 -7902 850 -7875
rect 899 -7902 916 -7875
rect -25 -7973 -8 -7946
rect 41 -7973 58 -7946
rect 107 -7973 124 -7946
rect 173 -7973 190 -7946
rect 239 -7973 256 -7946
rect 305 -7973 322 -7946
rect 371 -7973 388 -7946
rect 437 -7973 454 -7946
rect 503 -7973 520 -7946
rect 569 -7973 586 -7946
rect 635 -7973 652 -7946
rect 701 -7973 718 -7946
rect 767 -7973 784 -7946
rect 833 -7973 850 -7946
rect 899 -7973 916 -7946
rect -25 -8044 -8 -8017
rect 41 -8044 58 -8017
rect 107 -8044 124 -8017
rect 173 -8044 190 -8017
rect 239 -8044 256 -8017
rect 305 -8044 322 -8017
rect 371 -8044 388 -8017
rect 437 -8044 454 -8017
rect 503 -8044 520 -8017
rect 569 -8044 586 -8017
rect 635 -8044 652 -8017
rect 701 -8044 718 -8017
rect 767 -8044 784 -8017
rect 833 -8044 850 -8017
rect 899 -8044 916 -8017
rect -25 -8115 -8 -8088
rect 41 -8115 58 -8088
rect 107 -8115 124 -8088
rect 173 -8115 190 -8088
rect 239 -8115 256 -8088
rect 305 -8115 322 -8088
rect 371 -8115 388 -8088
rect 437 -8115 454 -8088
rect 503 -8115 520 -8088
rect 569 -8115 586 -8088
rect 635 -8115 652 -8088
rect 701 -8115 718 -8088
rect 767 -8115 784 -8088
rect 833 -8115 850 -8088
rect 899 -8115 916 -8088
rect -25 -8186 -8 -8159
rect 41 -8186 58 -8159
rect 107 -8186 124 -8159
rect 173 -8186 190 -8159
rect 239 -8186 256 -8159
rect 305 -8186 322 -8159
rect 371 -8186 388 -8159
rect 437 -8186 454 -8159
rect 503 -8186 520 -8159
rect 569 -8186 586 -8159
rect 635 -8186 652 -8159
rect 701 -8186 718 -8159
rect 767 -8186 784 -8159
rect 833 -8186 850 -8159
rect 899 -8186 916 -8159
rect -25 -8257 -8 -8230
rect 41 -8257 58 -8230
rect 107 -8257 124 -8230
rect 173 -8257 190 -8230
rect 239 -8257 256 -8230
rect 305 -8257 322 -8230
rect 371 -8257 388 -8230
rect 437 -8257 454 -8230
rect 503 -8257 520 -8230
rect 569 -8257 586 -8230
rect 635 -8257 652 -8230
rect 701 -8257 718 -8230
rect 767 -8257 784 -8230
rect 833 -8257 850 -8230
rect 899 -8257 916 -8230
rect -25 -8328 -8 -8301
rect 41 -8328 58 -8301
rect 107 -8328 124 -8301
rect 173 -8328 190 -8301
rect 239 -8328 256 -8301
rect 305 -8328 322 -8301
rect 371 -8328 388 -8301
rect 437 -8328 454 -8301
rect 503 -8328 520 -8301
rect 569 -8328 586 -8301
rect 635 -8328 652 -8301
rect 701 -8328 718 -8301
rect 767 -8328 784 -8301
rect 833 -8328 850 -8301
rect 899 -8328 916 -8301
rect -25 -8399 -8 -8372
rect 41 -8399 58 -8372
rect 107 -8399 124 -8372
rect 173 -8399 190 -8372
rect 239 -8399 256 -8372
rect 305 -8399 322 -8372
rect 371 -8399 388 -8372
rect 437 -8399 454 -8372
rect 503 -8399 520 -8372
rect 569 -8399 586 -8372
rect 635 -8399 652 -8372
rect 701 -8399 718 -8372
rect 767 -8399 784 -8372
rect 833 -8399 850 -8372
rect 899 -8399 916 -8372
rect -25 -8470 -8 -8443
rect 41 -8470 58 -8443
rect 107 -8470 124 -8443
rect 173 -8470 190 -8443
rect 239 -8470 256 -8443
rect 305 -8470 322 -8443
rect 371 -8470 388 -8443
rect 437 -8470 454 -8443
rect 503 -8470 520 -8443
rect 569 -8470 586 -8443
rect 635 -8470 652 -8443
rect 701 -8470 718 -8443
rect 767 -8470 784 -8443
rect 833 -8470 850 -8443
rect 899 -8470 916 -8443
rect -25 -8541 -8 -8514
rect 41 -8541 58 -8514
rect 107 -8541 124 -8514
rect 173 -8541 190 -8514
rect 239 -8541 256 -8514
rect 305 -8541 322 -8514
rect 371 -8541 388 -8514
rect 437 -8541 454 -8514
rect 503 -8541 520 -8514
rect 569 -8541 586 -8514
rect 635 -8541 652 -8514
rect 701 -8541 718 -8514
rect 767 -8541 784 -8514
rect 833 -8541 850 -8514
rect 899 -8541 916 -8514
rect -25 -8612 -8 -8585
rect 41 -8612 58 -8585
rect 107 -8612 124 -8585
rect 173 -8612 190 -8585
rect 239 -8612 256 -8585
rect 305 -8612 322 -8585
rect 371 -8612 388 -8585
rect 437 -8612 454 -8585
rect 503 -8612 520 -8585
rect 569 -8612 586 -8585
rect 635 -8612 652 -8585
rect 701 -8612 718 -8585
rect 767 -8612 784 -8585
rect 833 -8612 850 -8585
rect 899 -8612 916 -8585
rect -25 -8683 -8 -8656
rect 41 -8683 58 -8656
rect 107 -8683 124 -8656
rect 173 -8683 190 -8656
rect 239 -8683 256 -8656
rect 305 -8683 322 -8656
rect 371 -8683 388 -8656
rect 437 -8683 454 -8656
rect 503 -8683 520 -8656
rect 569 -8683 586 -8656
rect 635 -8683 652 -8656
rect 701 -8683 718 -8656
rect 767 -8683 784 -8656
rect 833 -8683 850 -8656
rect 899 -8683 916 -8656
rect -25 -8754 -8 -8727
rect 41 -8754 58 -8727
rect 107 -8754 124 -8727
rect 173 -8754 190 -8727
rect 239 -8754 256 -8727
rect 305 -8754 322 -8727
rect 371 -8754 388 -8727
rect 437 -8754 454 -8727
rect 503 -8754 520 -8727
rect 569 -8754 586 -8727
rect 635 -8754 652 -8727
rect 701 -8754 718 -8727
rect 767 -8754 784 -8727
rect 833 -8754 850 -8727
rect 899 -8754 916 -8727
rect -25 -8825 -8 -8798
rect 41 -8825 58 -8798
rect 107 -8825 124 -8798
rect 173 -8825 190 -8798
rect 239 -8825 256 -8798
rect 305 -8825 322 -8798
rect 371 -8825 388 -8798
rect 437 -8825 454 -8798
rect 503 -8825 520 -8798
rect 569 -8825 586 -8798
rect 635 -8825 652 -8798
rect 701 -8825 718 -8798
rect 767 -8825 784 -8798
rect 833 -8825 850 -8798
rect 899 -8825 916 -8798
rect -25 -8896 -8 -8869
rect 41 -8896 58 -8869
rect 107 -8896 124 -8869
rect 173 -8896 190 -8869
rect 239 -8896 256 -8869
rect 305 -8896 322 -8869
rect 371 -8896 388 -8869
rect 437 -8896 454 -8869
rect 503 -8896 520 -8869
rect 569 -8896 586 -8869
rect 635 -8896 652 -8869
rect 701 -8896 718 -8869
rect 767 -8896 784 -8869
rect 833 -8896 850 -8869
rect 899 -8896 916 -8869
rect -25 -8967 -8 -8940
rect 41 -8967 58 -8940
rect 107 -8967 124 -8940
rect 173 -8967 190 -8940
rect 239 -8967 256 -8940
rect 305 -8967 322 -8940
rect 371 -8967 388 -8940
rect 437 -8967 454 -8940
rect 503 -8967 520 -8940
rect 569 -8967 586 -8940
rect 635 -8967 652 -8940
rect 701 -8967 718 -8940
rect 767 -8967 784 -8940
rect 833 -8967 850 -8940
rect 899 -8967 916 -8940
rect -25 -9038 -8 -9011
rect 41 -9038 58 -9011
rect 107 -9038 124 -9011
rect 173 -9038 190 -9011
rect 239 -9038 256 -9011
rect 305 -9038 322 -9011
rect 371 -9038 388 -9011
rect 437 -9038 454 -9011
rect 503 -9038 520 -9011
rect 569 -9038 586 -9011
rect 635 -9038 652 -9011
rect 701 -9038 718 -9011
rect 767 -9038 784 -9011
rect 833 -9038 850 -9011
rect 899 -9038 916 -9011
rect -25 -9109 -8 -9082
rect 41 -9109 58 -9082
rect 107 -9109 124 -9082
rect 173 -9109 190 -9082
rect 239 -9109 256 -9082
rect 305 -9109 322 -9082
rect 371 -9109 388 -9082
rect 437 -9109 454 -9082
rect 503 -9109 520 -9082
rect 569 -9109 586 -9082
rect 635 -9109 652 -9082
rect 701 -9109 718 -9082
rect 767 -9109 784 -9082
rect 833 -9109 850 -9082
rect 899 -9109 916 -9082
rect 64 90 81 117
rect 8 90 25 117
rect 196 90 213 117
rect 140 90 157 117
rect 328 90 345 117
rect 272 90 289 117
rect 460 90 477 117
rect 404 90 421 117
rect 592 90 609 117
rect 536 90 553 117
rect 724 90 741 117
rect 668 90 685 117
rect 856 90 873 117
rect 800 90 817 117
rect 1073 90 1090 117
rect 1129 90 1146 117
rect 1205 90 1222 117
rect 1261 90 1278 117
rect 1337 90 1354 117
rect 1393 90 1410 117
rect 1469 90 1486 117
rect 1525 90 1542 117
rect 1601 90 1618 117
rect 1657 90 1674 117
rect 1733 90 1750 117
rect 1789 90 1806 117
rect 1865 90 1882 117
rect 1921 90 1938 117
<< ndiffc >>
rect 1030 -92 1047 -65
rect 1096 -92 1113 -65
rect 1162 -92 1179 -65
rect 1228 -92 1245 -65
rect 1294 -92 1311 -65
rect 1360 -92 1377 -65
rect 1426 -92 1443 -65
rect 1492 -92 1509 -65
rect 1558 -92 1575 -65
rect 1624 -92 1641 -65
rect 1690 -92 1707 -65
rect 1756 -92 1773 -65
rect 1822 -92 1839 -65
rect 1888 -92 1905 -65
rect 1162 -163 1179 -136
rect 1096 -163 1113 -136
rect 1162 -163 1179 -136
rect 1228 -163 1245 -136
rect 1294 -163 1311 -136
rect 1360 -163 1377 -136
rect 1426 -163 1443 -136
rect 1492 -163 1509 -136
rect 1558 -163 1575 -136
rect 1624 -163 1641 -136
rect 1690 -163 1707 -136
rect 1756 -163 1773 -136
rect 1822 -163 1839 -136
rect 1888 -163 1905 -136
rect 1030 -234 1047 -207
rect 1096 -234 1113 -207
rect 1294 -234 1311 -207
rect 1228 -234 1245 -207
rect 1294 -234 1311 -207
rect 1360 -234 1377 -207
rect 1426 -234 1443 -207
rect 1492 -234 1509 -207
rect 1558 -234 1575 -207
rect 1624 -234 1641 -207
rect 1690 -234 1707 -207
rect 1756 -234 1773 -207
rect 1822 -234 1839 -207
rect 1888 -234 1905 -207
rect 1162 -305 1179 -278
rect 1096 -305 1113 -278
rect 1294 -305 1311 -278
rect 1228 -305 1245 -278
rect 1294 -305 1311 -278
rect 1360 -305 1377 -278
rect 1426 -305 1443 -278
rect 1492 -305 1509 -278
rect 1558 -305 1575 -278
rect 1624 -305 1641 -278
rect 1690 -305 1707 -278
rect 1756 -305 1773 -278
rect 1822 -305 1839 -278
rect 1888 -305 1905 -278
rect 1030 -376 1047 -349
rect 1096 -376 1113 -349
rect 1162 -376 1179 -349
rect 1228 -376 1245 -349
rect 1426 -376 1443 -349
rect 1360 -376 1377 -349
rect 1426 -376 1443 -349
rect 1492 -376 1509 -349
rect 1558 -376 1575 -349
rect 1624 -376 1641 -349
rect 1690 -376 1707 -349
rect 1756 -376 1773 -349
rect 1822 -376 1839 -349
rect 1888 -376 1905 -349
rect 1162 -447 1179 -420
rect 1096 -447 1113 -420
rect 1162 -447 1179 -420
rect 1228 -447 1245 -420
rect 1426 -447 1443 -420
rect 1360 -447 1377 -420
rect 1426 -447 1443 -420
rect 1492 -447 1509 -420
rect 1558 -447 1575 -420
rect 1624 -447 1641 -420
rect 1690 -447 1707 -420
rect 1756 -447 1773 -420
rect 1822 -447 1839 -420
rect 1888 -447 1905 -420
rect 1030 -518 1047 -491
rect 1096 -518 1113 -491
rect 1294 -518 1311 -491
rect 1228 -518 1245 -491
rect 1426 -518 1443 -491
rect 1360 -518 1377 -491
rect 1426 -518 1443 -491
rect 1492 -518 1509 -491
rect 1558 -518 1575 -491
rect 1624 -518 1641 -491
rect 1690 -518 1707 -491
rect 1756 -518 1773 -491
rect 1822 -518 1839 -491
rect 1888 -518 1905 -491
rect 1162 -589 1179 -562
rect 1096 -589 1113 -562
rect 1294 -589 1311 -562
rect 1228 -589 1245 -562
rect 1426 -589 1443 -562
rect 1360 -589 1377 -562
rect 1426 -589 1443 -562
rect 1492 -589 1509 -562
rect 1558 -589 1575 -562
rect 1624 -589 1641 -562
rect 1690 -589 1707 -562
rect 1756 -589 1773 -562
rect 1822 -589 1839 -562
rect 1888 -589 1905 -562
rect 1030 -660 1047 -633
rect 1096 -660 1113 -633
rect 1162 -660 1179 -633
rect 1228 -660 1245 -633
rect 1294 -660 1311 -633
rect 1360 -660 1377 -633
rect 1558 -660 1575 -633
rect 1492 -660 1509 -633
rect 1558 -660 1575 -633
rect 1624 -660 1641 -633
rect 1690 -660 1707 -633
rect 1756 -660 1773 -633
rect 1822 -660 1839 -633
rect 1888 -660 1905 -633
rect 1162 -731 1179 -704
rect 1096 -731 1113 -704
rect 1162 -731 1179 -704
rect 1228 -731 1245 -704
rect 1294 -731 1311 -704
rect 1360 -731 1377 -704
rect 1558 -731 1575 -704
rect 1492 -731 1509 -704
rect 1558 -731 1575 -704
rect 1624 -731 1641 -704
rect 1690 -731 1707 -704
rect 1756 -731 1773 -704
rect 1822 -731 1839 -704
rect 1888 -731 1905 -704
rect 1030 -802 1047 -775
rect 1096 -802 1113 -775
rect 1294 -802 1311 -775
rect 1228 -802 1245 -775
rect 1294 -802 1311 -775
rect 1360 -802 1377 -775
rect 1558 -802 1575 -775
rect 1492 -802 1509 -775
rect 1558 -802 1575 -775
rect 1624 -802 1641 -775
rect 1690 -802 1707 -775
rect 1756 -802 1773 -775
rect 1822 -802 1839 -775
rect 1888 -802 1905 -775
rect 1162 -873 1179 -846
rect 1096 -873 1113 -846
rect 1294 -873 1311 -846
rect 1228 -873 1245 -846
rect 1294 -873 1311 -846
rect 1360 -873 1377 -846
rect 1558 -873 1575 -846
rect 1492 -873 1509 -846
rect 1558 -873 1575 -846
rect 1624 -873 1641 -846
rect 1690 -873 1707 -846
rect 1756 -873 1773 -846
rect 1822 -873 1839 -846
rect 1888 -873 1905 -846
rect 1030 -944 1047 -917
rect 1096 -944 1113 -917
rect 1162 -944 1179 -917
rect 1228 -944 1245 -917
rect 1426 -944 1443 -917
rect 1360 -944 1377 -917
rect 1558 -944 1575 -917
rect 1492 -944 1509 -917
rect 1558 -944 1575 -917
rect 1624 -944 1641 -917
rect 1690 -944 1707 -917
rect 1756 -944 1773 -917
rect 1822 -944 1839 -917
rect 1888 -944 1905 -917
rect 1162 -1015 1179 -988
rect 1096 -1015 1113 -988
rect 1162 -1015 1179 -988
rect 1228 -1015 1245 -988
rect 1426 -1015 1443 -988
rect 1360 -1015 1377 -988
rect 1558 -1015 1575 -988
rect 1492 -1015 1509 -988
rect 1558 -1015 1575 -988
rect 1624 -1015 1641 -988
rect 1690 -1015 1707 -988
rect 1756 -1015 1773 -988
rect 1822 -1015 1839 -988
rect 1888 -1015 1905 -988
rect 1030 -1086 1047 -1059
rect 1096 -1086 1113 -1059
rect 1294 -1086 1311 -1059
rect 1228 -1086 1245 -1059
rect 1426 -1086 1443 -1059
rect 1360 -1086 1377 -1059
rect 1558 -1086 1575 -1059
rect 1492 -1086 1509 -1059
rect 1558 -1086 1575 -1059
rect 1624 -1086 1641 -1059
rect 1690 -1086 1707 -1059
rect 1756 -1086 1773 -1059
rect 1822 -1086 1839 -1059
rect 1888 -1086 1905 -1059
rect 1162 -1157 1179 -1130
rect 1096 -1157 1113 -1130
rect 1294 -1157 1311 -1130
rect 1228 -1157 1245 -1130
rect 1426 -1157 1443 -1130
rect 1360 -1157 1377 -1130
rect 1558 -1157 1575 -1130
rect 1492 -1157 1509 -1130
rect 1558 -1157 1575 -1130
rect 1624 -1157 1641 -1130
rect 1690 -1157 1707 -1130
rect 1756 -1157 1773 -1130
rect 1822 -1157 1839 -1130
rect 1888 -1157 1905 -1130
rect 1030 -1228 1047 -1201
rect 1096 -1228 1113 -1201
rect 1162 -1228 1179 -1201
rect 1228 -1228 1245 -1201
rect 1294 -1228 1311 -1201
rect 1360 -1228 1377 -1201
rect 1426 -1228 1443 -1201
rect 1492 -1228 1509 -1201
rect 1690 -1228 1707 -1201
rect 1624 -1228 1641 -1201
rect 1690 -1228 1707 -1201
rect 1756 -1228 1773 -1201
rect 1822 -1228 1839 -1201
rect 1888 -1228 1905 -1201
rect 1162 -1299 1179 -1272
rect 1096 -1299 1113 -1272
rect 1162 -1299 1179 -1272
rect 1228 -1299 1245 -1272
rect 1294 -1299 1311 -1272
rect 1360 -1299 1377 -1272
rect 1426 -1299 1443 -1272
rect 1492 -1299 1509 -1272
rect 1690 -1299 1707 -1272
rect 1624 -1299 1641 -1272
rect 1690 -1299 1707 -1272
rect 1756 -1299 1773 -1272
rect 1822 -1299 1839 -1272
rect 1888 -1299 1905 -1272
rect 1030 -1370 1047 -1343
rect 1096 -1370 1113 -1343
rect 1294 -1370 1311 -1343
rect 1228 -1370 1245 -1343
rect 1294 -1370 1311 -1343
rect 1360 -1370 1377 -1343
rect 1426 -1370 1443 -1343
rect 1492 -1370 1509 -1343
rect 1690 -1370 1707 -1343
rect 1624 -1370 1641 -1343
rect 1690 -1370 1707 -1343
rect 1756 -1370 1773 -1343
rect 1822 -1370 1839 -1343
rect 1888 -1370 1905 -1343
rect 1162 -1441 1179 -1414
rect 1096 -1441 1113 -1414
rect 1294 -1441 1311 -1414
rect 1228 -1441 1245 -1414
rect 1294 -1441 1311 -1414
rect 1360 -1441 1377 -1414
rect 1426 -1441 1443 -1414
rect 1492 -1441 1509 -1414
rect 1690 -1441 1707 -1414
rect 1624 -1441 1641 -1414
rect 1690 -1441 1707 -1414
rect 1756 -1441 1773 -1414
rect 1822 -1441 1839 -1414
rect 1888 -1441 1905 -1414
rect 1030 -1512 1047 -1485
rect 1096 -1512 1113 -1485
rect 1162 -1512 1179 -1485
rect 1228 -1512 1245 -1485
rect 1426 -1512 1443 -1485
rect 1360 -1512 1377 -1485
rect 1426 -1512 1443 -1485
rect 1492 -1512 1509 -1485
rect 1690 -1512 1707 -1485
rect 1624 -1512 1641 -1485
rect 1690 -1512 1707 -1485
rect 1756 -1512 1773 -1485
rect 1822 -1512 1839 -1485
rect 1888 -1512 1905 -1485
rect 1162 -1583 1179 -1556
rect 1096 -1583 1113 -1556
rect 1162 -1583 1179 -1556
rect 1228 -1583 1245 -1556
rect 1426 -1583 1443 -1556
rect 1360 -1583 1377 -1556
rect 1426 -1583 1443 -1556
rect 1492 -1583 1509 -1556
rect 1690 -1583 1707 -1556
rect 1624 -1583 1641 -1556
rect 1690 -1583 1707 -1556
rect 1756 -1583 1773 -1556
rect 1822 -1583 1839 -1556
rect 1888 -1583 1905 -1556
rect 1030 -1654 1047 -1627
rect 1096 -1654 1113 -1627
rect 1294 -1654 1311 -1627
rect 1228 -1654 1245 -1627
rect 1426 -1654 1443 -1627
rect 1360 -1654 1377 -1627
rect 1426 -1654 1443 -1627
rect 1492 -1654 1509 -1627
rect 1690 -1654 1707 -1627
rect 1624 -1654 1641 -1627
rect 1690 -1654 1707 -1627
rect 1756 -1654 1773 -1627
rect 1822 -1654 1839 -1627
rect 1888 -1654 1905 -1627
rect 1162 -1725 1179 -1698
rect 1096 -1725 1113 -1698
rect 1294 -1725 1311 -1698
rect 1228 -1725 1245 -1698
rect 1426 -1725 1443 -1698
rect 1360 -1725 1377 -1698
rect 1426 -1725 1443 -1698
rect 1492 -1725 1509 -1698
rect 1690 -1725 1707 -1698
rect 1624 -1725 1641 -1698
rect 1690 -1725 1707 -1698
rect 1756 -1725 1773 -1698
rect 1822 -1725 1839 -1698
rect 1888 -1725 1905 -1698
rect 1030 -1796 1047 -1769
rect 1096 -1796 1113 -1769
rect 1162 -1796 1179 -1769
rect 1228 -1796 1245 -1769
rect 1294 -1796 1311 -1769
rect 1360 -1796 1377 -1769
rect 1558 -1796 1575 -1769
rect 1492 -1796 1509 -1769
rect 1690 -1796 1707 -1769
rect 1624 -1796 1641 -1769
rect 1690 -1796 1707 -1769
rect 1756 -1796 1773 -1769
rect 1822 -1796 1839 -1769
rect 1888 -1796 1905 -1769
rect 1162 -1867 1179 -1840
rect 1096 -1867 1113 -1840
rect 1162 -1867 1179 -1840
rect 1228 -1867 1245 -1840
rect 1294 -1867 1311 -1840
rect 1360 -1867 1377 -1840
rect 1558 -1867 1575 -1840
rect 1492 -1867 1509 -1840
rect 1690 -1867 1707 -1840
rect 1624 -1867 1641 -1840
rect 1690 -1867 1707 -1840
rect 1756 -1867 1773 -1840
rect 1822 -1867 1839 -1840
rect 1888 -1867 1905 -1840
rect 1030 -1938 1047 -1911
rect 1096 -1938 1113 -1911
rect 1294 -1938 1311 -1911
rect 1228 -1938 1245 -1911
rect 1294 -1938 1311 -1911
rect 1360 -1938 1377 -1911
rect 1558 -1938 1575 -1911
rect 1492 -1938 1509 -1911
rect 1690 -1938 1707 -1911
rect 1624 -1938 1641 -1911
rect 1690 -1938 1707 -1911
rect 1756 -1938 1773 -1911
rect 1822 -1938 1839 -1911
rect 1888 -1938 1905 -1911
rect 1162 -2009 1179 -1982
rect 1096 -2009 1113 -1982
rect 1294 -2009 1311 -1982
rect 1228 -2009 1245 -1982
rect 1294 -2009 1311 -1982
rect 1360 -2009 1377 -1982
rect 1558 -2009 1575 -1982
rect 1492 -2009 1509 -1982
rect 1690 -2009 1707 -1982
rect 1624 -2009 1641 -1982
rect 1690 -2009 1707 -1982
rect 1756 -2009 1773 -1982
rect 1822 -2009 1839 -1982
rect 1888 -2009 1905 -1982
rect 1030 -2080 1047 -2053
rect 1096 -2080 1113 -2053
rect 1162 -2080 1179 -2053
rect 1228 -2080 1245 -2053
rect 1426 -2080 1443 -2053
rect 1360 -2080 1377 -2053
rect 1558 -2080 1575 -2053
rect 1492 -2080 1509 -2053
rect 1690 -2080 1707 -2053
rect 1624 -2080 1641 -2053
rect 1690 -2080 1707 -2053
rect 1756 -2080 1773 -2053
rect 1822 -2080 1839 -2053
rect 1888 -2080 1905 -2053
rect 1162 -2151 1179 -2124
rect 1096 -2151 1113 -2124
rect 1162 -2151 1179 -2124
rect 1228 -2151 1245 -2124
rect 1426 -2151 1443 -2124
rect 1360 -2151 1377 -2124
rect 1558 -2151 1575 -2124
rect 1492 -2151 1509 -2124
rect 1690 -2151 1707 -2124
rect 1624 -2151 1641 -2124
rect 1690 -2151 1707 -2124
rect 1756 -2151 1773 -2124
rect 1822 -2151 1839 -2124
rect 1888 -2151 1905 -2124
rect 1030 -2222 1047 -2195
rect 1096 -2222 1113 -2195
rect 1294 -2222 1311 -2195
rect 1228 -2222 1245 -2195
rect 1426 -2222 1443 -2195
rect 1360 -2222 1377 -2195
rect 1558 -2222 1575 -2195
rect 1492 -2222 1509 -2195
rect 1690 -2222 1707 -2195
rect 1624 -2222 1641 -2195
rect 1690 -2222 1707 -2195
rect 1756 -2222 1773 -2195
rect 1822 -2222 1839 -2195
rect 1888 -2222 1905 -2195
rect 1162 -2293 1179 -2266
rect 1096 -2293 1113 -2266
rect 1294 -2293 1311 -2266
rect 1228 -2293 1245 -2266
rect 1426 -2293 1443 -2266
rect 1360 -2293 1377 -2266
rect 1558 -2293 1575 -2266
rect 1492 -2293 1509 -2266
rect 1690 -2293 1707 -2266
rect 1624 -2293 1641 -2266
rect 1690 -2293 1707 -2266
rect 1756 -2293 1773 -2266
rect 1822 -2293 1839 -2266
rect 1888 -2293 1905 -2266
rect 1030 -2364 1047 -2337
rect 1096 -2364 1113 -2337
rect 1162 -2364 1179 -2337
rect 1228 -2364 1245 -2337
rect 1294 -2364 1311 -2337
rect 1360 -2364 1377 -2337
rect 1426 -2364 1443 -2337
rect 1492 -2364 1509 -2337
rect 1558 -2364 1575 -2337
rect 1624 -2364 1641 -2337
rect 1822 -2364 1839 -2337
rect 1756 -2364 1773 -2337
rect 1822 -2364 1839 -2337
rect 1888 -2364 1905 -2337
rect 1162 -2435 1179 -2408
rect 1096 -2435 1113 -2408
rect 1162 -2435 1179 -2408
rect 1228 -2435 1245 -2408
rect 1294 -2435 1311 -2408
rect 1360 -2435 1377 -2408
rect 1426 -2435 1443 -2408
rect 1492 -2435 1509 -2408
rect 1558 -2435 1575 -2408
rect 1624 -2435 1641 -2408
rect 1822 -2435 1839 -2408
rect 1756 -2435 1773 -2408
rect 1822 -2435 1839 -2408
rect 1888 -2435 1905 -2408
rect 1030 -2506 1047 -2479
rect 1096 -2506 1113 -2479
rect 1294 -2506 1311 -2479
rect 1228 -2506 1245 -2479
rect 1294 -2506 1311 -2479
rect 1360 -2506 1377 -2479
rect 1426 -2506 1443 -2479
rect 1492 -2506 1509 -2479
rect 1558 -2506 1575 -2479
rect 1624 -2506 1641 -2479
rect 1822 -2506 1839 -2479
rect 1756 -2506 1773 -2479
rect 1822 -2506 1839 -2479
rect 1888 -2506 1905 -2479
rect 1162 -2577 1179 -2550
rect 1096 -2577 1113 -2550
rect 1294 -2577 1311 -2550
rect 1228 -2577 1245 -2550
rect 1294 -2577 1311 -2550
rect 1360 -2577 1377 -2550
rect 1426 -2577 1443 -2550
rect 1492 -2577 1509 -2550
rect 1558 -2577 1575 -2550
rect 1624 -2577 1641 -2550
rect 1822 -2577 1839 -2550
rect 1756 -2577 1773 -2550
rect 1822 -2577 1839 -2550
rect 1888 -2577 1905 -2550
rect 1030 -2648 1047 -2621
rect 1096 -2648 1113 -2621
rect 1162 -2648 1179 -2621
rect 1228 -2648 1245 -2621
rect 1426 -2648 1443 -2621
rect 1360 -2648 1377 -2621
rect 1426 -2648 1443 -2621
rect 1492 -2648 1509 -2621
rect 1558 -2648 1575 -2621
rect 1624 -2648 1641 -2621
rect 1822 -2648 1839 -2621
rect 1756 -2648 1773 -2621
rect 1822 -2648 1839 -2621
rect 1888 -2648 1905 -2621
rect 1162 -2719 1179 -2692
rect 1096 -2719 1113 -2692
rect 1162 -2719 1179 -2692
rect 1228 -2719 1245 -2692
rect 1426 -2719 1443 -2692
rect 1360 -2719 1377 -2692
rect 1426 -2719 1443 -2692
rect 1492 -2719 1509 -2692
rect 1558 -2719 1575 -2692
rect 1624 -2719 1641 -2692
rect 1822 -2719 1839 -2692
rect 1756 -2719 1773 -2692
rect 1822 -2719 1839 -2692
rect 1888 -2719 1905 -2692
rect 1030 -2790 1047 -2763
rect 1096 -2790 1113 -2763
rect 1294 -2790 1311 -2763
rect 1228 -2790 1245 -2763
rect 1426 -2790 1443 -2763
rect 1360 -2790 1377 -2763
rect 1426 -2790 1443 -2763
rect 1492 -2790 1509 -2763
rect 1558 -2790 1575 -2763
rect 1624 -2790 1641 -2763
rect 1822 -2790 1839 -2763
rect 1756 -2790 1773 -2763
rect 1822 -2790 1839 -2763
rect 1888 -2790 1905 -2763
rect 1162 -2861 1179 -2834
rect 1096 -2861 1113 -2834
rect 1294 -2861 1311 -2834
rect 1228 -2861 1245 -2834
rect 1426 -2861 1443 -2834
rect 1360 -2861 1377 -2834
rect 1426 -2861 1443 -2834
rect 1492 -2861 1509 -2834
rect 1558 -2861 1575 -2834
rect 1624 -2861 1641 -2834
rect 1822 -2861 1839 -2834
rect 1756 -2861 1773 -2834
rect 1822 -2861 1839 -2834
rect 1888 -2861 1905 -2834
rect 1030 -2932 1047 -2905
rect 1096 -2932 1113 -2905
rect 1162 -2932 1179 -2905
rect 1228 -2932 1245 -2905
rect 1294 -2932 1311 -2905
rect 1360 -2932 1377 -2905
rect 1558 -2932 1575 -2905
rect 1492 -2932 1509 -2905
rect 1558 -2932 1575 -2905
rect 1624 -2932 1641 -2905
rect 1822 -2932 1839 -2905
rect 1756 -2932 1773 -2905
rect 1822 -2932 1839 -2905
rect 1888 -2932 1905 -2905
rect 1162 -3003 1179 -2976
rect 1096 -3003 1113 -2976
rect 1162 -3003 1179 -2976
rect 1228 -3003 1245 -2976
rect 1294 -3003 1311 -2976
rect 1360 -3003 1377 -2976
rect 1558 -3003 1575 -2976
rect 1492 -3003 1509 -2976
rect 1558 -3003 1575 -2976
rect 1624 -3003 1641 -2976
rect 1822 -3003 1839 -2976
rect 1756 -3003 1773 -2976
rect 1822 -3003 1839 -2976
rect 1888 -3003 1905 -2976
rect 1030 -3074 1047 -3047
rect 1096 -3074 1113 -3047
rect 1294 -3074 1311 -3047
rect 1228 -3074 1245 -3047
rect 1294 -3074 1311 -3047
rect 1360 -3074 1377 -3047
rect 1558 -3074 1575 -3047
rect 1492 -3074 1509 -3047
rect 1558 -3074 1575 -3047
rect 1624 -3074 1641 -3047
rect 1822 -3074 1839 -3047
rect 1756 -3074 1773 -3047
rect 1822 -3074 1839 -3047
rect 1888 -3074 1905 -3047
rect 1162 -3145 1179 -3118
rect 1096 -3145 1113 -3118
rect 1294 -3145 1311 -3118
rect 1228 -3145 1245 -3118
rect 1294 -3145 1311 -3118
rect 1360 -3145 1377 -3118
rect 1558 -3145 1575 -3118
rect 1492 -3145 1509 -3118
rect 1558 -3145 1575 -3118
rect 1624 -3145 1641 -3118
rect 1822 -3145 1839 -3118
rect 1756 -3145 1773 -3118
rect 1822 -3145 1839 -3118
rect 1888 -3145 1905 -3118
rect 1030 -3216 1047 -3189
rect 1096 -3216 1113 -3189
rect 1162 -3216 1179 -3189
rect 1228 -3216 1245 -3189
rect 1426 -3216 1443 -3189
rect 1360 -3216 1377 -3189
rect 1558 -3216 1575 -3189
rect 1492 -3216 1509 -3189
rect 1558 -3216 1575 -3189
rect 1624 -3216 1641 -3189
rect 1822 -3216 1839 -3189
rect 1756 -3216 1773 -3189
rect 1822 -3216 1839 -3189
rect 1888 -3216 1905 -3189
rect 1162 -3287 1179 -3260
rect 1096 -3287 1113 -3260
rect 1162 -3287 1179 -3260
rect 1228 -3287 1245 -3260
rect 1426 -3287 1443 -3260
rect 1360 -3287 1377 -3260
rect 1558 -3287 1575 -3260
rect 1492 -3287 1509 -3260
rect 1558 -3287 1575 -3260
rect 1624 -3287 1641 -3260
rect 1822 -3287 1839 -3260
rect 1756 -3287 1773 -3260
rect 1822 -3287 1839 -3260
rect 1888 -3287 1905 -3260
rect 1030 -3358 1047 -3331
rect 1096 -3358 1113 -3331
rect 1294 -3358 1311 -3331
rect 1228 -3358 1245 -3331
rect 1426 -3358 1443 -3331
rect 1360 -3358 1377 -3331
rect 1558 -3358 1575 -3331
rect 1492 -3358 1509 -3331
rect 1558 -3358 1575 -3331
rect 1624 -3358 1641 -3331
rect 1822 -3358 1839 -3331
rect 1756 -3358 1773 -3331
rect 1822 -3358 1839 -3331
rect 1888 -3358 1905 -3331
rect 1162 -3429 1179 -3402
rect 1096 -3429 1113 -3402
rect 1294 -3429 1311 -3402
rect 1228 -3429 1245 -3402
rect 1426 -3429 1443 -3402
rect 1360 -3429 1377 -3402
rect 1558 -3429 1575 -3402
rect 1492 -3429 1509 -3402
rect 1558 -3429 1575 -3402
rect 1624 -3429 1641 -3402
rect 1822 -3429 1839 -3402
rect 1756 -3429 1773 -3402
rect 1822 -3429 1839 -3402
rect 1888 -3429 1905 -3402
rect 1030 -3500 1047 -3473
rect 1096 -3500 1113 -3473
rect 1162 -3500 1179 -3473
rect 1228 -3500 1245 -3473
rect 1294 -3500 1311 -3473
rect 1360 -3500 1377 -3473
rect 1426 -3500 1443 -3473
rect 1492 -3500 1509 -3473
rect 1690 -3500 1707 -3473
rect 1624 -3500 1641 -3473
rect 1822 -3500 1839 -3473
rect 1756 -3500 1773 -3473
rect 1822 -3500 1839 -3473
rect 1888 -3500 1905 -3473
rect 1162 -3571 1179 -3544
rect 1096 -3571 1113 -3544
rect 1162 -3571 1179 -3544
rect 1228 -3571 1245 -3544
rect 1294 -3571 1311 -3544
rect 1360 -3571 1377 -3544
rect 1426 -3571 1443 -3544
rect 1492 -3571 1509 -3544
rect 1690 -3571 1707 -3544
rect 1624 -3571 1641 -3544
rect 1822 -3571 1839 -3544
rect 1756 -3571 1773 -3544
rect 1822 -3571 1839 -3544
rect 1888 -3571 1905 -3544
rect 1030 -3642 1047 -3615
rect 1096 -3642 1113 -3615
rect 1294 -3642 1311 -3615
rect 1228 -3642 1245 -3615
rect 1294 -3642 1311 -3615
rect 1360 -3642 1377 -3615
rect 1426 -3642 1443 -3615
rect 1492 -3642 1509 -3615
rect 1690 -3642 1707 -3615
rect 1624 -3642 1641 -3615
rect 1822 -3642 1839 -3615
rect 1756 -3642 1773 -3615
rect 1822 -3642 1839 -3615
rect 1888 -3642 1905 -3615
rect 1162 -3713 1179 -3686
rect 1096 -3713 1113 -3686
rect 1294 -3713 1311 -3686
rect 1228 -3713 1245 -3686
rect 1294 -3713 1311 -3686
rect 1360 -3713 1377 -3686
rect 1426 -3713 1443 -3686
rect 1492 -3713 1509 -3686
rect 1690 -3713 1707 -3686
rect 1624 -3713 1641 -3686
rect 1822 -3713 1839 -3686
rect 1756 -3713 1773 -3686
rect 1822 -3713 1839 -3686
rect 1888 -3713 1905 -3686
rect 1030 -3784 1047 -3757
rect 1096 -3784 1113 -3757
rect 1162 -3784 1179 -3757
rect 1228 -3784 1245 -3757
rect 1426 -3784 1443 -3757
rect 1360 -3784 1377 -3757
rect 1426 -3784 1443 -3757
rect 1492 -3784 1509 -3757
rect 1690 -3784 1707 -3757
rect 1624 -3784 1641 -3757
rect 1822 -3784 1839 -3757
rect 1756 -3784 1773 -3757
rect 1822 -3784 1839 -3757
rect 1888 -3784 1905 -3757
rect 1162 -3855 1179 -3828
rect 1096 -3855 1113 -3828
rect 1162 -3855 1179 -3828
rect 1228 -3855 1245 -3828
rect 1426 -3855 1443 -3828
rect 1360 -3855 1377 -3828
rect 1426 -3855 1443 -3828
rect 1492 -3855 1509 -3828
rect 1690 -3855 1707 -3828
rect 1624 -3855 1641 -3828
rect 1822 -3855 1839 -3828
rect 1756 -3855 1773 -3828
rect 1822 -3855 1839 -3828
rect 1888 -3855 1905 -3828
rect 1030 -3926 1047 -3899
rect 1096 -3926 1113 -3899
rect 1294 -3926 1311 -3899
rect 1228 -3926 1245 -3899
rect 1426 -3926 1443 -3899
rect 1360 -3926 1377 -3899
rect 1426 -3926 1443 -3899
rect 1492 -3926 1509 -3899
rect 1690 -3926 1707 -3899
rect 1624 -3926 1641 -3899
rect 1822 -3926 1839 -3899
rect 1756 -3926 1773 -3899
rect 1822 -3926 1839 -3899
rect 1888 -3926 1905 -3899
rect 1162 -3997 1179 -3970
rect 1096 -3997 1113 -3970
rect 1294 -3997 1311 -3970
rect 1228 -3997 1245 -3970
rect 1426 -3997 1443 -3970
rect 1360 -3997 1377 -3970
rect 1426 -3997 1443 -3970
rect 1492 -3997 1509 -3970
rect 1690 -3997 1707 -3970
rect 1624 -3997 1641 -3970
rect 1822 -3997 1839 -3970
rect 1756 -3997 1773 -3970
rect 1822 -3997 1839 -3970
rect 1888 -3997 1905 -3970
rect 1030 -4068 1047 -4041
rect 1096 -4068 1113 -4041
rect 1162 -4068 1179 -4041
rect 1228 -4068 1245 -4041
rect 1294 -4068 1311 -4041
rect 1360 -4068 1377 -4041
rect 1558 -4068 1575 -4041
rect 1492 -4068 1509 -4041
rect 1690 -4068 1707 -4041
rect 1624 -4068 1641 -4041
rect 1822 -4068 1839 -4041
rect 1756 -4068 1773 -4041
rect 1822 -4068 1839 -4041
rect 1888 -4068 1905 -4041
rect 1162 -4139 1179 -4112
rect 1096 -4139 1113 -4112
rect 1162 -4139 1179 -4112
rect 1228 -4139 1245 -4112
rect 1294 -4139 1311 -4112
rect 1360 -4139 1377 -4112
rect 1558 -4139 1575 -4112
rect 1492 -4139 1509 -4112
rect 1690 -4139 1707 -4112
rect 1624 -4139 1641 -4112
rect 1822 -4139 1839 -4112
rect 1756 -4139 1773 -4112
rect 1822 -4139 1839 -4112
rect 1888 -4139 1905 -4112
rect 1030 -4210 1047 -4183
rect 1096 -4210 1113 -4183
rect 1294 -4210 1311 -4183
rect 1228 -4210 1245 -4183
rect 1294 -4210 1311 -4183
rect 1360 -4210 1377 -4183
rect 1558 -4210 1575 -4183
rect 1492 -4210 1509 -4183
rect 1690 -4210 1707 -4183
rect 1624 -4210 1641 -4183
rect 1822 -4210 1839 -4183
rect 1756 -4210 1773 -4183
rect 1822 -4210 1839 -4183
rect 1888 -4210 1905 -4183
rect 1162 -4281 1179 -4254
rect 1096 -4281 1113 -4254
rect 1294 -4281 1311 -4254
rect 1228 -4281 1245 -4254
rect 1294 -4281 1311 -4254
rect 1360 -4281 1377 -4254
rect 1558 -4281 1575 -4254
rect 1492 -4281 1509 -4254
rect 1690 -4281 1707 -4254
rect 1624 -4281 1641 -4254
rect 1822 -4281 1839 -4254
rect 1756 -4281 1773 -4254
rect 1822 -4281 1839 -4254
rect 1888 -4281 1905 -4254
rect 1030 -4352 1047 -4325
rect 1096 -4352 1113 -4325
rect 1162 -4352 1179 -4325
rect 1228 -4352 1245 -4325
rect 1426 -4352 1443 -4325
rect 1360 -4352 1377 -4325
rect 1558 -4352 1575 -4325
rect 1492 -4352 1509 -4325
rect 1690 -4352 1707 -4325
rect 1624 -4352 1641 -4325
rect 1822 -4352 1839 -4325
rect 1756 -4352 1773 -4325
rect 1822 -4352 1839 -4325
rect 1888 -4352 1905 -4325
rect 1162 -4423 1179 -4396
rect 1096 -4423 1113 -4396
rect 1162 -4423 1179 -4396
rect 1228 -4423 1245 -4396
rect 1426 -4423 1443 -4396
rect 1360 -4423 1377 -4396
rect 1558 -4423 1575 -4396
rect 1492 -4423 1509 -4396
rect 1690 -4423 1707 -4396
rect 1624 -4423 1641 -4396
rect 1822 -4423 1839 -4396
rect 1756 -4423 1773 -4396
rect 1822 -4423 1839 -4396
rect 1888 -4423 1905 -4396
rect 1030 -4494 1047 -4467
rect 1096 -4494 1113 -4467
rect 1294 -4494 1311 -4467
rect 1228 -4494 1245 -4467
rect 1426 -4494 1443 -4467
rect 1360 -4494 1377 -4467
rect 1558 -4494 1575 -4467
rect 1492 -4494 1509 -4467
rect 1690 -4494 1707 -4467
rect 1624 -4494 1641 -4467
rect 1822 -4494 1839 -4467
rect 1756 -4494 1773 -4467
rect 1822 -4494 1839 -4467
rect 1888 -4494 1905 -4467
rect 1162 -4565 1179 -4538
rect 1096 -4565 1113 -4538
rect 1294 -4565 1311 -4538
rect 1228 -4565 1245 -4538
rect 1426 -4565 1443 -4538
rect 1360 -4565 1377 -4538
rect 1558 -4565 1575 -4538
rect 1492 -4565 1509 -4538
rect 1690 -4565 1707 -4538
rect 1624 -4565 1641 -4538
rect 1822 -4565 1839 -4538
rect 1756 -4565 1773 -4538
rect 1822 -4565 1839 -4538
rect 1888 -4565 1905 -4538
rect 1030 -4636 1047 -4609
rect 1096 -4636 1113 -4609
rect 1162 -4636 1179 -4609
rect 1228 -4636 1245 -4609
rect 1294 -4636 1311 -4609
rect 1360 -4636 1377 -4609
rect 1426 -4636 1443 -4609
rect 1492 -4636 1509 -4609
rect 1558 -4636 1575 -4609
rect 1624 -4636 1641 -4609
rect 1690 -4636 1707 -4609
rect 1756 -4636 1773 -4609
rect 1954 -4636 1971 -4609
rect 1954 -4636 1971 -4609
rect 1888 -4636 1905 -4609
rect 1162 -4707 1179 -4680
rect 1096 -4707 1113 -4680
rect 1162 -4707 1179 -4680
rect 1228 -4707 1245 -4680
rect 1294 -4707 1311 -4680
rect 1360 -4707 1377 -4680
rect 1426 -4707 1443 -4680
rect 1492 -4707 1509 -4680
rect 1558 -4707 1575 -4680
rect 1624 -4707 1641 -4680
rect 1690 -4707 1707 -4680
rect 1756 -4707 1773 -4680
rect 1954 -4707 1971 -4680
rect 1954 -4707 1971 -4680
rect 1888 -4707 1905 -4680
rect 1030 -4778 1047 -4751
rect 1096 -4778 1113 -4751
rect 1294 -4778 1311 -4751
rect 1228 -4778 1245 -4751
rect 1294 -4778 1311 -4751
rect 1360 -4778 1377 -4751
rect 1426 -4778 1443 -4751
rect 1492 -4778 1509 -4751
rect 1558 -4778 1575 -4751
rect 1624 -4778 1641 -4751
rect 1690 -4778 1707 -4751
rect 1756 -4778 1773 -4751
rect 1954 -4778 1971 -4751
rect 1954 -4778 1971 -4751
rect 1888 -4778 1905 -4751
rect 1162 -4849 1179 -4822
rect 1096 -4849 1113 -4822
rect 1294 -4849 1311 -4822
rect 1228 -4849 1245 -4822
rect 1294 -4849 1311 -4822
rect 1360 -4849 1377 -4822
rect 1426 -4849 1443 -4822
rect 1492 -4849 1509 -4822
rect 1558 -4849 1575 -4822
rect 1624 -4849 1641 -4822
rect 1690 -4849 1707 -4822
rect 1756 -4849 1773 -4822
rect 1954 -4849 1971 -4822
rect 1954 -4849 1971 -4822
rect 1888 -4849 1905 -4822
rect 1030 -4920 1047 -4893
rect 1096 -4920 1113 -4893
rect 1162 -4920 1179 -4893
rect 1228 -4920 1245 -4893
rect 1426 -4920 1443 -4893
rect 1360 -4920 1377 -4893
rect 1426 -4920 1443 -4893
rect 1492 -4920 1509 -4893
rect 1558 -4920 1575 -4893
rect 1624 -4920 1641 -4893
rect 1690 -4920 1707 -4893
rect 1756 -4920 1773 -4893
rect 1954 -4920 1971 -4893
rect 1954 -4920 1971 -4893
rect 1888 -4920 1905 -4893
rect 1162 -4991 1179 -4964
rect 1096 -4991 1113 -4964
rect 1162 -4991 1179 -4964
rect 1228 -4991 1245 -4964
rect 1426 -4991 1443 -4964
rect 1360 -4991 1377 -4964
rect 1426 -4991 1443 -4964
rect 1492 -4991 1509 -4964
rect 1558 -4991 1575 -4964
rect 1624 -4991 1641 -4964
rect 1690 -4991 1707 -4964
rect 1756 -4991 1773 -4964
rect 1954 -4991 1971 -4964
rect 1954 -4991 1971 -4964
rect 1888 -4991 1905 -4964
rect 1030 -5062 1047 -5035
rect 1096 -5062 1113 -5035
rect 1294 -5062 1311 -5035
rect 1228 -5062 1245 -5035
rect 1426 -5062 1443 -5035
rect 1360 -5062 1377 -5035
rect 1426 -5062 1443 -5035
rect 1492 -5062 1509 -5035
rect 1558 -5062 1575 -5035
rect 1624 -5062 1641 -5035
rect 1690 -5062 1707 -5035
rect 1756 -5062 1773 -5035
rect 1954 -5062 1971 -5035
rect 1954 -5062 1971 -5035
rect 1888 -5062 1905 -5035
rect 1162 -5133 1179 -5106
rect 1096 -5133 1113 -5106
rect 1294 -5133 1311 -5106
rect 1228 -5133 1245 -5106
rect 1426 -5133 1443 -5106
rect 1360 -5133 1377 -5106
rect 1426 -5133 1443 -5106
rect 1492 -5133 1509 -5106
rect 1558 -5133 1575 -5106
rect 1624 -5133 1641 -5106
rect 1690 -5133 1707 -5106
rect 1756 -5133 1773 -5106
rect 1954 -5133 1971 -5106
rect 1954 -5133 1971 -5106
rect 1888 -5133 1905 -5106
rect 1030 -5204 1047 -5177
rect 1096 -5204 1113 -5177
rect 1162 -5204 1179 -5177
rect 1228 -5204 1245 -5177
rect 1294 -5204 1311 -5177
rect 1360 -5204 1377 -5177
rect 1558 -5204 1575 -5177
rect 1492 -5204 1509 -5177
rect 1558 -5204 1575 -5177
rect 1624 -5204 1641 -5177
rect 1690 -5204 1707 -5177
rect 1756 -5204 1773 -5177
rect 1954 -5204 1971 -5177
rect 1954 -5204 1971 -5177
rect 1888 -5204 1905 -5177
rect 1162 -5275 1179 -5248
rect 1096 -5275 1113 -5248
rect 1162 -5275 1179 -5248
rect 1228 -5275 1245 -5248
rect 1294 -5275 1311 -5248
rect 1360 -5275 1377 -5248
rect 1558 -5275 1575 -5248
rect 1492 -5275 1509 -5248
rect 1558 -5275 1575 -5248
rect 1624 -5275 1641 -5248
rect 1690 -5275 1707 -5248
rect 1756 -5275 1773 -5248
rect 1954 -5275 1971 -5248
rect 1954 -5275 1971 -5248
rect 1888 -5275 1905 -5248
rect 1030 -5346 1047 -5319
rect 1096 -5346 1113 -5319
rect 1294 -5346 1311 -5319
rect 1228 -5346 1245 -5319
rect 1294 -5346 1311 -5319
rect 1360 -5346 1377 -5319
rect 1558 -5346 1575 -5319
rect 1492 -5346 1509 -5319
rect 1558 -5346 1575 -5319
rect 1624 -5346 1641 -5319
rect 1690 -5346 1707 -5319
rect 1756 -5346 1773 -5319
rect 1954 -5346 1971 -5319
rect 1954 -5346 1971 -5319
rect 1888 -5346 1905 -5319
rect 1162 -5417 1179 -5390
rect 1096 -5417 1113 -5390
rect 1294 -5417 1311 -5390
rect 1228 -5417 1245 -5390
rect 1294 -5417 1311 -5390
rect 1360 -5417 1377 -5390
rect 1558 -5417 1575 -5390
rect 1492 -5417 1509 -5390
rect 1558 -5417 1575 -5390
rect 1624 -5417 1641 -5390
rect 1690 -5417 1707 -5390
rect 1756 -5417 1773 -5390
rect 1954 -5417 1971 -5390
rect 1954 -5417 1971 -5390
rect 1888 -5417 1905 -5390
rect 1030 -5488 1047 -5461
rect 1096 -5488 1113 -5461
rect 1162 -5488 1179 -5461
rect 1228 -5488 1245 -5461
rect 1426 -5488 1443 -5461
rect 1360 -5488 1377 -5461
rect 1558 -5488 1575 -5461
rect 1492 -5488 1509 -5461
rect 1558 -5488 1575 -5461
rect 1624 -5488 1641 -5461
rect 1690 -5488 1707 -5461
rect 1756 -5488 1773 -5461
rect 1954 -5488 1971 -5461
rect 1954 -5488 1971 -5461
rect 1888 -5488 1905 -5461
rect 1162 -5559 1179 -5532
rect 1096 -5559 1113 -5532
rect 1162 -5559 1179 -5532
rect 1228 -5559 1245 -5532
rect 1426 -5559 1443 -5532
rect 1360 -5559 1377 -5532
rect 1558 -5559 1575 -5532
rect 1492 -5559 1509 -5532
rect 1558 -5559 1575 -5532
rect 1624 -5559 1641 -5532
rect 1690 -5559 1707 -5532
rect 1756 -5559 1773 -5532
rect 1954 -5559 1971 -5532
rect 1954 -5559 1971 -5532
rect 1888 -5559 1905 -5532
rect 1030 -5630 1047 -5603
rect 1096 -5630 1113 -5603
rect 1294 -5630 1311 -5603
rect 1228 -5630 1245 -5603
rect 1426 -5630 1443 -5603
rect 1360 -5630 1377 -5603
rect 1558 -5630 1575 -5603
rect 1492 -5630 1509 -5603
rect 1558 -5630 1575 -5603
rect 1624 -5630 1641 -5603
rect 1690 -5630 1707 -5603
rect 1756 -5630 1773 -5603
rect 1954 -5630 1971 -5603
rect 1954 -5630 1971 -5603
rect 1888 -5630 1905 -5603
rect 1162 -5701 1179 -5674
rect 1096 -5701 1113 -5674
rect 1294 -5701 1311 -5674
rect 1228 -5701 1245 -5674
rect 1426 -5701 1443 -5674
rect 1360 -5701 1377 -5674
rect 1558 -5701 1575 -5674
rect 1492 -5701 1509 -5674
rect 1558 -5701 1575 -5674
rect 1624 -5701 1641 -5674
rect 1690 -5701 1707 -5674
rect 1756 -5701 1773 -5674
rect 1954 -5701 1971 -5674
rect 1954 -5701 1971 -5674
rect 1888 -5701 1905 -5674
rect 1030 -5772 1047 -5745
rect 1096 -5772 1113 -5745
rect 1162 -5772 1179 -5745
rect 1228 -5772 1245 -5745
rect 1294 -5772 1311 -5745
rect 1360 -5772 1377 -5745
rect 1426 -5772 1443 -5745
rect 1492 -5772 1509 -5745
rect 1690 -5772 1707 -5745
rect 1624 -5772 1641 -5745
rect 1690 -5772 1707 -5745
rect 1756 -5772 1773 -5745
rect 1954 -5772 1971 -5745
rect 1954 -5772 1971 -5745
rect 1888 -5772 1905 -5745
rect 1162 -5843 1179 -5816
rect 1096 -5843 1113 -5816
rect 1162 -5843 1179 -5816
rect 1228 -5843 1245 -5816
rect 1294 -5843 1311 -5816
rect 1360 -5843 1377 -5816
rect 1426 -5843 1443 -5816
rect 1492 -5843 1509 -5816
rect 1690 -5843 1707 -5816
rect 1624 -5843 1641 -5816
rect 1690 -5843 1707 -5816
rect 1756 -5843 1773 -5816
rect 1954 -5843 1971 -5816
rect 1954 -5843 1971 -5816
rect 1888 -5843 1905 -5816
rect 1030 -5914 1047 -5887
rect 1096 -5914 1113 -5887
rect 1294 -5914 1311 -5887
rect 1228 -5914 1245 -5887
rect 1294 -5914 1311 -5887
rect 1360 -5914 1377 -5887
rect 1426 -5914 1443 -5887
rect 1492 -5914 1509 -5887
rect 1690 -5914 1707 -5887
rect 1624 -5914 1641 -5887
rect 1690 -5914 1707 -5887
rect 1756 -5914 1773 -5887
rect 1954 -5914 1971 -5887
rect 1954 -5914 1971 -5887
rect 1888 -5914 1905 -5887
rect 1162 -5985 1179 -5958
rect 1096 -5985 1113 -5958
rect 1294 -5985 1311 -5958
rect 1228 -5985 1245 -5958
rect 1294 -5985 1311 -5958
rect 1360 -5985 1377 -5958
rect 1426 -5985 1443 -5958
rect 1492 -5985 1509 -5958
rect 1690 -5985 1707 -5958
rect 1624 -5985 1641 -5958
rect 1690 -5985 1707 -5958
rect 1756 -5985 1773 -5958
rect 1954 -5985 1971 -5958
rect 1954 -5985 1971 -5958
rect 1888 -5985 1905 -5958
rect 1030 -6056 1047 -6029
rect 1096 -6056 1113 -6029
rect 1162 -6056 1179 -6029
rect 1228 -6056 1245 -6029
rect 1426 -6056 1443 -6029
rect 1360 -6056 1377 -6029
rect 1426 -6056 1443 -6029
rect 1492 -6056 1509 -6029
rect 1690 -6056 1707 -6029
rect 1624 -6056 1641 -6029
rect 1690 -6056 1707 -6029
rect 1756 -6056 1773 -6029
rect 1954 -6056 1971 -6029
rect 1954 -6056 1971 -6029
rect 1888 -6056 1905 -6029
rect 1162 -6127 1179 -6100
rect 1096 -6127 1113 -6100
rect 1162 -6127 1179 -6100
rect 1228 -6127 1245 -6100
rect 1426 -6127 1443 -6100
rect 1360 -6127 1377 -6100
rect 1426 -6127 1443 -6100
rect 1492 -6127 1509 -6100
rect 1690 -6127 1707 -6100
rect 1624 -6127 1641 -6100
rect 1690 -6127 1707 -6100
rect 1756 -6127 1773 -6100
rect 1954 -6127 1971 -6100
rect 1954 -6127 1971 -6100
rect 1888 -6127 1905 -6100
rect 1030 -6198 1047 -6171
rect 1096 -6198 1113 -6171
rect 1294 -6198 1311 -6171
rect 1228 -6198 1245 -6171
rect 1426 -6198 1443 -6171
rect 1360 -6198 1377 -6171
rect 1426 -6198 1443 -6171
rect 1492 -6198 1509 -6171
rect 1690 -6198 1707 -6171
rect 1624 -6198 1641 -6171
rect 1690 -6198 1707 -6171
rect 1756 -6198 1773 -6171
rect 1954 -6198 1971 -6171
rect 1954 -6198 1971 -6171
rect 1888 -6198 1905 -6171
rect 1162 -6269 1179 -6242
rect 1096 -6269 1113 -6242
rect 1294 -6269 1311 -6242
rect 1228 -6269 1245 -6242
rect 1426 -6269 1443 -6242
rect 1360 -6269 1377 -6242
rect 1426 -6269 1443 -6242
rect 1492 -6269 1509 -6242
rect 1690 -6269 1707 -6242
rect 1624 -6269 1641 -6242
rect 1690 -6269 1707 -6242
rect 1756 -6269 1773 -6242
rect 1954 -6269 1971 -6242
rect 1954 -6269 1971 -6242
rect 1888 -6269 1905 -6242
rect 1030 -6340 1047 -6313
rect 1096 -6340 1113 -6313
rect 1162 -6340 1179 -6313
rect 1228 -6340 1245 -6313
rect 1294 -6340 1311 -6313
rect 1360 -6340 1377 -6313
rect 1558 -6340 1575 -6313
rect 1492 -6340 1509 -6313
rect 1690 -6340 1707 -6313
rect 1624 -6340 1641 -6313
rect 1690 -6340 1707 -6313
rect 1756 -6340 1773 -6313
rect 1954 -6340 1971 -6313
rect 1954 -6340 1971 -6313
rect 1888 -6340 1905 -6313
rect 1162 -6411 1179 -6384
rect 1096 -6411 1113 -6384
rect 1162 -6411 1179 -6384
rect 1228 -6411 1245 -6384
rect 1294 -6411 1311 -6384
rect 1360 -6411 1377 -6384
rect 1558 -6411 1575 -6384
rect 1492 -6411 1509 -6384
rect 1690 -6411 1707 -6384
rect 1624 -6411 1641 -6384
rect 1690 -6411 1707 -6384
rect 1756 -6411 1773 -6384
rect 1954 -6411 1971 -6384
rect 1954 -6411 1971 -6384
rect 1888 -6411 1905 -6384
rect 1030 -6482 1047 -6455
rect 1096 -6482 1113 -6455
rect 1294 -6482 1311 -6455
rect 1228 -6482 1245 -6455
rect 1294 -6482 1311 -6455
rect 1360 -6482 1377 -6455
rect 1558 -6482 1575 -6455
rect 1492 -6482 1509 -6455
rect 1690 -6482 1707 -6455
rect 1624 -6482 1641 -6455
rect 1690 -6482 1707 -6455
rect 1756 -6482 1773 -6455
rect 1954 -6482 1971 -6455
rect 1954 -6482 1971 -6455
rect 1888 -6482 1905 -6455
rect 1162 -6553 1179 -6526
rect 1096 -6553 1113 -6526
rect 1294 -6553 1311 -6526
rect 1228 -6553 1245 -6526
rect 1294 -6553 1311 -6526
rect 1360 -6553 1377 -6526
rect 1558 -6553 1575 -6526
rect 1492 -6553 1509 -6526
rect 1690 -6553 1707 -6526
rect 1624 -6553 1641 -6526
rect 1690 -6553 1707 -6526
rect 1756 -6553 1773 -6526
rect 1954 -6553 1971 -6526
rect 1954 -6553 1971 -6526
rect 1888 -6553 1905 -6526
rect 1030 -6624 1047 -6597
rect 1096 -6624 1113 -6597
rect 1162 -6624 1179 -6597
rect 1228 -6624 1245 -6597
rect 1426 -6624 1443 -6597
rect 1360 -6624 1377 -6597
rect 1558 -6624 1575 -6597
rect 1492 -6624 1509 -6597
rect 1690 -6624 1707 -6597
rect 1624 -6624 1641 -6597
rect 1690 -6624 1707 -6597
rect 1756 -6624 1773 -6597
rect 1954 -6624 1971 -6597
rect 1954 -6624 1971 -6597
rect 1888 -6624 1905 -6597
rect 1162 -6695 1179 -6668
rect 1096 -6695 1113 -6668
rect 1162 -6695 1179 -6668
rect 1228 -6695 1245 -6668
rect 1426 -6695 1443 -6668
rect 1360 -6695 1377 -6668
rect 1558 -6695 1575 -6668
rect 1492 -6695 1509 -6668
rect 1690 -6695 1707 -6668
rect 1624 -6695 1641 -6668
rect 1690 -6695 1707 -6668
rect 1756 -6695 1773 -6668
rect 1954 -6695 1971 -6668
rect 1954 -6695 1971 -6668
rect 1888 -6695 1905 -6668
rect 1030 -6766 1047 -6739
rect 1096 -6766 1113 -6739
rect 1294 -6766 1311 -6739
rect 1228 -6766 1245 -6739
rect 1426 -6766 1443 -6739
rect 1360 -6766 1377 -6739
rect 1558 -6766 1575 -6739
rect 1492 -6766 1509 -6739
rect 1690 -6766 1707 -6739
rect 1624 -6766 1641 -6739
rect 1690 -6766 1707 -6739
rect 1756 -6766 1773 -6739
rect 1954 -6766 1971 -6739
rect 1954 -6766 1971 -6739
rect 1888 -6766 1905 -6739
rect 1162 -6837 1179 -6810
rect 1096 -6837 1113 -6810
rect 1294 -6837 1311 -6810
rect 1228 -6837 1245 -6810
rect 1426 -6837 1443 -6810
rect 1360 -6837 1377 -6810
rect 1558 -6837 1575 -6810
rect 1492 -6837 1509 -6810
rect 1690 -6837 1707 -6810
rect 1624 -6837 1641 -6810
rect 1690 -6837 1707 -6810
rect 1756 -6837 1773 -6810
rect 1954 -6837 1971 -6810
rect 1954 -6837 1971 -6810
rect 1888 -6837 1905 -6810
rect 1030 -6908 1047 -6881
rect 1096 -6908 1113 -6881
rect 1162 -6908 1179 -6881
rect 1228 -6908 1245 -6881
rect 1294 -6908 1311 -6881
rect 1360 -6908 1377 -6881
rect 1426 -6908 1443 -6881
rect 1492 -6908 1509 -6881
rect 1558 -6908 1575 -6881
rect 1624 -6908 1641 -6881
rect 1822 -6908 1839 -6881
rect 1756 -6908 1773 -6881
rect 1954 -6908 1971 -6881
rect 1954 -6908 1971 -6881
rect 1888 -6908 1905 -6881
rect 1162 -6979 1179 -6952
rect 1096 -6979 1113 -6952
rect 1162 -6979 1179 -6952
rect 1228 -6979 1245 -6952
rect 1294 -6979 1311 -6952
rect 1360 -6979 1377 -6952
rect 1426 -6979 1443 -6952
rect 1492 -6979 1509 -6952
rect 1558 -6979 1575 -6952
rect 1624 -6979 1641 -6952
rect 1822 -6979 1839 -6952
rect 1756 -6979 1773 -6952
rect 1954 -6979 1971 -6952
rect 1954 -6979 1971 -6952
rect 1888 -6979 1905 -6952
rect 1030 -7050 1047 -7023
rect 1096 -7050 1113 -7023
rect 1294 -7050 1311 -7023
rect 1228 -7050 1245 -7023
rect 1294 -7050 1311 -7023
rect 1360 -7050 1377 -7023
rect 1426 -7050 1443 -7023
rect 1492 -7050 1509 -7023
rect 1558 -7050 1575 -7023
rect 1624 -7050 1641 -7023
rect 1822 -7050 1839 -7023
rect 1756 -7050 1773 -7023
rect 1954 -7050 1971 -7023
rect 1954 -7050 1971 -7023
rect 1888 -7050 1905 -7023
rect 1162 -7121 1179 -7094
rect 1096 -7121 1113 -7094
rect 1294 -7121 1311 -7094
rect 1228 -7121 1245 -7094
rect 1294 -7121 1311 -7094
rect 1360 -7121 1377 -7094
rect 1426 -7121 1443 -7094
rect 1492 -7121 1509 -7094
rect 1558 -7121 1575 -7094
rect 1624 -7121 1641 -7094
rect 1822 -7121 1839 -7094
rect 1756 -7121 1773 -7094
rect 1954 -7121 1971 -7094
rect 1954 -7121 1971 -7094
rect 1888 -7121 1905 -7094
rect 1030 -7192 1047 -7165
rect 1096 -7192 1113 -7165
rect 1162 -7192 1179 -7165
rect 1228 -7192 1245 -7165
rect 1426 -7192 1443 -7165
rect 1360 -7192 1377 -7165
rect 1426 -7192 1443 -7165
rect 1492 -7192 1509 -7165
rect 1558 -7192 1575 -7165
rect 1624 -7192 1641 -7165
rect 1822 -7192 1839 -7165
rect 1756 -7192 1773 -7165
rect 1954 -7192 1971 -7165
rect 1954 -7192 1971 -7165
rect 1888 -7192 1905 -7165
rect 1162 -7263 1179 -7236
rect 1096 -7263 1113 -7236
rect 1162 -7263 1179 -7236
rect 1228 -7263 1245 -7236
rect 1426 -7263 1443 -7236
rect 1360 -7263 1377 -7236
rect 1426 -7263 1443 -7236
rect 1492 -7263 1509 -7236
rect 1558 -7263 1575 -7236
rect 1624 -7263 1641 -7236
rect 1822 -7263 1839 -7236
rect 1756 -7263 1773 -7236
rect 1954 -7263 1971 -7236
rect 1954 -7263 1971 -7236
rect 1888 -7263 1905 -7236
rect 1030 -7334 1047 -7307
rect 1096 -7334 1113 -7307
rect 1294 -7334 1311 -7307
rect 1228 -7334 1245 -7307
rect 1426 -7334 1443 -7307
rect 1360 -7334 1377 -7307
rect 1426 -7334 1443 -7307
rect 1492 -7334 1509 -7307
rect 1558 -7334 1575 -7307
rect 1624 -7334 1641 -7307
rect 1822 -7334 1839 -7307
rect 1756 -7334 1773 -7307
rect 1954 -7334 1971 -7307
rect 1954 -7334 1971 -7307
rect 1888 -7334 1905 -7307
rect 1162 -7405 1179 -7378
rect 1096 -7405 1113 -7378
rect 1294 -7405 1311 -7378
rect 1228 -7405 1245 -7378
rect 1426 -7405 1443 -7378
rect 1360 -7405 1377 -7378
rect 1426 -7405 1443 -7378
rect 1492 -7405 1509 -7378
rect 1558 -7405 1575 -7378
rect 1624 -7405 1641 -7378
rect 1822 -7405 1839 -7378
rect 1756 -7405 1773 -7378
rect 1954 -7405 1971 -7378
rect 1954 -7405 1971 -7378
rect 1888 -7405 1905 -7378
rect 1030 -7476 1047 -7449
rect 1096 -7476 1113 -7449
rect 1162 -7476 1179 -7449
rect 1228 -7476 1245 -7449
rect 1294 -7476 1311 -7449
rect 1360 -7476 1377 -7449
rect 1558 -7476 1575 -7449
rect 1492 -7476 1509 -7449
rect 1558 -7476 1575 -7449
rect 1624 -7476 1641 -7449
rect 1822 -7476 1839 -7449
rect 1756 -7476 1773 -7449
rect 1954 -7476 1971 -7449
rect 1954 -7476 1971 -7449
rect 1888 -7476 1905 -7449
rect 1162 -7547 1179 -7520
rect 1096 -7547 1113 -7520
rect 1162 -7547 1179 -7520
rect 1228 -7547 1245 -7520
rect 1294 -7547 1311 -7520
rect 1360 -7547 1377 -7520
rect 1558 -7547 1575 -7520
rect 1492 -7547 1509 -7520
rect 1558 -7547 1575 -7520
rect 1624 -7547 1641 -7520
rect 1822 -7547 1839 -7520
rect 1756 -7547 1773 -7520
rect 1954 -7547 1971 -7520
rect 1954 -7547 1971 -7520
rect 1888 -7547 1905 -7520
rect 1030 -7618 1047 -7591
rect 1096 -7618 1113 -7591
rect 1294 -7618 1311 -7591
rect 1228 -7618 1245 -7591
rect 1294 -7618 1311 -7591
rect 1360 -7618 1377 -7591
rect 1558 -7618 1575 -7591
rect 1492 -7618 1509 -7591
rect 1558 -7618 1575 -7591
rect 1624 -7618 1641 -7591
rect 1822 -7618 1839 -7591
rect 1756 -7618 1773 -7591
rect 1954 -7618 1971 -7591
rect 1954 -7618 1971 -7591
rect 1888 -7618 1905 -7591
rect 1162 -7689 1179 -7662
rect 1096 -7689 1113 -7662
rect 1294 -7689 1311 -7662
rect 1228 -7689 1245 -7662
rect 1294 -7689 1311 -7662
rect 1360 -7689 1377 -7662
rect 1558 -7689 1575 -7662
rect 1492 -7689 1509 -7662
rect 1558 -7689 1575 -7662
rect 1624 -7689 1641 -7662
rect 1822 -7689 1839 -7662
rect 1756 -7689 1773 -7662
rect 1954 -7689 1971 -7662
rect 1954 -7689 1971 -7662
rect 1888 -7689 1905 -7662
rect 1030 -7760 1047 -7733
rect 1096 -7760 1113 -7733
rect 1162 -7760 1179 -7733
rect 1228 -7760 1245 -7733
rect 1426 -7760 1443 -7733
rect 1360 -7760 1377 -7733
rect 1558 -7760 1575 -7733
rect 1492 -7760 1509 -7733
rect 1558 -7760 1575 -7733
rect 1624 -7760 1641 -7733
rect 1822 -7760 1839 -7733
rect 1756 -7760 1773 -7733
rect 1954 -7760 1971 -7733
rect 1954 -7760 1971 -7733
rect 1888 -7760 1905 -7733
rect 1162 -7831 1179 -7804
rect 1096 -7831 1113 -7804
rect 1162 -7831 1179 -7804
rect 1228 -7831 1245 -7804
rect 1426 -7831 1443 -7804
rect 1360 -7831 1377 -7804
rect 1558 -7831 1575 -7804
rect 1492 -7831 1509 -7804
rect 1558 -7831 1575 -7804
rect 1624 -7831 1641 -7804
rect 1822 -7831 1839 -7804
rect 1756 -7831 1773 -7804
rect 1954 -7831 1971 -7804
rect 1954 -7831 1971 -7804
rect 1888 -7831 1905 -7804
rect 1030 -7902 1047 -7875
rect 1096 -7902 1113 -7875
rect 1294 -7902 1311 -7875
rect 1228 -7902 1245 -7875
rect 1426 -7902 1443 -7875
rect 1360 -7902 1377 -7875
rect 1558 -7902 1575 -7875
rect 1492 -7902 1509 -7875
rect 1558 -7902 1575 -7875
rect 1624 -7902 1641 -7875
rect 1822 -7902 1839 -7875
rect 1756 -7902 1773 -7875
rect 1954 -7902 1971 -7875
rect 1954 -7902 1971 -7875
rect 1888 -7902 1905 -7875
rect 1162 -7973 1179 -7946
rect 1096 -7973 1113 -7946
rect 1294 -7973 1311 -7946
rect 1228 -7973 1245 -7946
rect 1426 -7973 1443 -7946
rect 1360 -7973 1377 -7946
rect 1558 -7973 1575 -7946
rect 1492 -7973 1509 -7946
rect 1558 -7973 1575 -7946
rect 1624 -7973 1641 -7946
rect 1822 -7973 1839 -7946
rect 1756 -7973 1773 -7946
rect 1954 -7973 1971 -7946
rect 1954 -7973 1971 -7946
rect 1888 -7973 1905 -7946
rect 1030 -8044 1047 -8017
rect 1096 -8044 1113 -8017
rect 1162 -8044 1179 -8017
rect 1228 -8044 1245 -8017
rect 1294 -8044 1311 -8017
rect 1360 -8044 1377 -8017
rect 1426 -8044 1443 -8017
rect 1492 -8044 1509 -8017
rect 1690 -8044 1707 -8017
rect 1624 -8044 1641 -8017
rect 1822 -8044 1839 -8017
rect 1756 -8044 1773 -8017
rect 1954 -8044 1971 -8017
rect 1954 -8044 1971 -8017
rect 1888 -8044 1905 -8017
rect 1162 -8115 1179 -8088
rect 1096 -8115 1113 -8088
rect 1162 -8115 1179 -8088
rect 1228 -8115 1245 -8088
rect 1294 -8115 1311 -8088
rect 1360 -8115 1377 -8088
rect 1426 -8115 1443 -8088
rect 1492 -8115 1509 -8088
rect 1690 -8115 1707 -8088
rect 1624 -8115 1641 -8088
rect 1822 -8115 1839 -8088
rect 1756 -8115 1773 -8088
rect 1954 -8115 1971 -8088
rect 1954 -8115 1971 -8088
rect 1888 -8115 1905 -8088
rect 1030 -8186 1047 -8159
rect 1096 -8186 1113 -8159
rect 1294 -8186 1311 -8159
rect 1228 -8186 1245 -8159
rect 1294 -8186 1311 -8159
rect 1360 -8186 1377 -8159
rect 1426 -8186 1443 -8159
rect 1492 -8186 1509 -8159
rect 1690 -8186 1707 -8159
rect 1624 -8186 1641 -8159
rect 1822 -8186 1839 -8159
rect 1756 -8186 1773 -8159
rect 1954 -8186 1971 -8159
rect 1954 -8186 1971 -8159
rect 1888 -8186 1905 -8159
rect 1162 -8257 1179 -8230
rect 1096 -8257 1113 -8230
rect 1294 -8257 1311 -8230
rect 1228 -8257 1245 -8230
rect 1294 -8257 1311 -8230
rect 1360 -8257 1377 -8230
rect 1426 -8257 1443 -8230
rect 1492 -8257 1509 -8230
rect 1690 -8257 1707 -8230
rect 1624 -8257 1641 -8230
rect 1822 -8257 1839 -8230
rect 1756 -8257 1773 -8230
rect 1954 -8257 1971 -8230
rect 1954 -8257 1971 -8230
rect 1888 -8257 1905 -8230
rect 1030 -8328 1047 -8301
rect 1096 -8328 1113 -8301
rect 1162 -8328 1179 -8301
rect 1228 -8328 1245 -8301
rect 1426 -8328 1443 -8301
rect 1360 -8328 1377 -8301
rect 1426 -8328 1443 -8301
rect 1492 -8328 1509 -8301
rect 1690 -8328 1707 -8301
rect 1624 -8328 1641 -8301
rect 1822 -8328 1839 -8301
rect 1756 -8328 1773 -8301
rect 1954 -8328 1971 -8301
rect 1954 -8328 1971 -8301
rect 1888 -8328 1905 -8301
rect 1162 -8399 1179 -8372
rect 1096 -8399 1113 -8372
rect 1162 -8399 1179 -8372
rect 1228 -8399 1245 -8372
rect 1426 -8399 1443 -8372
rect 1360 -8399 1377 -8372
rect 1426 -8399 1443 -8372
rect 1492 -8399 1509 -8372
rect 1690 -8399 1707 -8372
rect 1624 -8399 1641 -8372
rect 1822 -8399 1839 -8372
rect 1756 -8399 1773 -8372
rect 1954 -8399 1971 -8372
rect 1954 -8399 1971 -8372
rect 1888 -8399 1905 -8372
rect 1030 -8470 1047 -8443
rect 1096 -8470 1113 -8443
rect 1294 -8470 1311 -8443
rect 1228 -8470 1245 -8443
rect 1426 -8470 1443 -8443
rect 1360 -8470 1377 -8443
rect 1426 -8470 1443 -8443
rect 1492 -8470 1509 -8443
rect 1690 -8470 1707 -8443
rect 1624 -8470 1641 -8443
rect 1822 -8470 1839 -8443
rect 1756 -8470 1773 -8443
rect 1954 -8470 1971 -8443
rect 1954 -8470 1971 -8443
rect 1888 -8470 1905 -8443
rect 1162 -8541 1179 -8514
rect 1096 -8541 1113 -8514
rect 1294 -8541 1311 -8514
rect 1228 -8541 1245 -8514
rect 1426 -8541 1443 -8514
rect 1360 -8541 1377 -8514
rect 1426 -8541 1443 -8514
rect 1492 -8541 1509 -8514
rect 1690 -8541 1707 -8514
rect 1624 -8541 1641 -8514
rect 1822 -8541 1839 -8514
rect 1756 -8541 1773 -8514
rect 1954 -8541 1971 -8514
rect 1954 -8541 1971 -8514
rect 1888 -8541 1905 -8514
rect 1030 -8612 1047 -8585
rect 1096 -8612 1113 -8585
rect 1162 -8612 1179 -8585
rect 1228 -8612 1245 -8585
rect 1294 -8612 1311 -8585
rect 1360 -8612 1377 -8585
rect 1558 -8612 1575 -8585
rect 1492 -8612 1509 -8585
rect 1690 -8612 1707 -8585
rect 1624 -8612 1641 -8585
rect 1822 -8612 1839 -8585
rect 1756 -8612 1773 -8585
rect 1954 -8612 1971 -8585
rect 1954 -8612 1971 -8585
rect 1888 -8612 1905 -8585
rect 1162 -8683 1179 -8656
rect 1096 -8683 1113 -8656
rect 1162 -8683 1179 -8656
rect 1228 -8683 1245 -8656
rect 1294 -8683 1311 -8656
rect 1360 -8683 1377 -8656
rect 1558 -8683 1575 -8656
rect 1492 -8683 1509 -8656
rect 1690 -8683 1707 -8656
rect 1624 -8683 1641 -8656
rect 1822 -8683 1839 -8656
rect 1756 -8683 1773 -8656
rect 1954 -8683 1971 -8656
rect 1954 -8683 1971 -8656
rect 1888 -8683 1905 -8656
rect 1030 -8754 1047 -8727
rect 1096 -8754 1113 -8727
rect 1294 -8754 1311 -8727
rect 1228 -8754 1245 -8727
rect 1294 -8754 1311 -8727
rect 1360 -8754 1377 -8727
rect 1558 -8754 1575 -8727
rect 1492 -8754 1509 -8727
rect 1690 -8754 1707 -8727
rect 1624 -8754 1641 -8727
rect 1822 -8754 1839 -8727
rect 1756 -8754 1773 -8727
rect 1954 -8754 1971 -8727
rect 1954 -8754 1971 -8727
rect 1888 -8754 1905 -8727
rect 1162 -8825 1179 -8798
rect 1096 -8825 1113 -8798
rect 1294 -8825 1311 -8798
rect 1228 -8825 1245 -8798
rect 1294 -8825 1311 -8798
rect 1360 -8825 1377 -8798
rect 1558 -8825 1575 -8798
rect 1492 -8825 1509 -8798
rect 1690 -8825 1707 -8798
rect 1624 -8825 1641 -8798
rect 1822 -8825 1839 -8798
rect 1756 -8825 1773 -8798
rect 1954 -8825 1971 -8798
rect 1954 -8825 1971 -8798
rect 1888 -8825 1905 -8798
rect 1030 -8896 1047 -8869
rect 1096 -8896 1113 -8869
rect 1162 -8896 1179 -8869
rect 1228 -8896 1245 -8869
rect 1426 -8896 1443 -8869
rect 1360 -8896 1377 -8869
rect 1558 -8896 1575 -8869
rect 1492 -8896 1509 -8869
rect 1690 -8896 1707 -8869
rect 1624 -8896 1641 -8869
rect 1822 -8896 1839 -8869
rect 1756 -8896 1773 -8869
rect 1954 -8896 1971 -8869
rect 1954 -8896 1971 -8869
rect 1888 -8896 1905 -8869
rect 1162 -8967 1179 -8940
rect 1096 -8967 1113 -8940
rect 1162 -8967 1179 -8940
rect 1228 -8967 1245 -8940
rect 1426 -8967 1443 -8940
rect 1360 -8967 1377 -8940
rect 1558 -8967 1575 -8940
rect 1492 -8967 1509 -8940
rect 1690 -8967 1707 -8940
rect 1624 -8967 1641 -8940
rect 1822 -8967 1839 -8940
rect 1756 -8967 1773 -8940
rect 1954 -8967 1971 -8940
rect 1954 -8967 1971 -8940
rect 1888 -8967 1905 -8940
rect 1030 -9038 1047 -9011
rect 1096 -9038 1113 -9011
rect 1294 -9038 1311 -9011
rect 1228 -9038 1245 -9011
rect 1426 -9038 1443 -9011
rect 1360 -9038 1377 -9011
rect 1558 -9038 1575 -9011
rect 1492 -9038 1509 -9011
rect 1690 -9038 1707 -9011
rect 1624 -9038 1641 -9011
rect 1822 -9038 1839 -9011
rect 1756 -9038 1773 -9011
rect 1954 -9038 1971 -9011
rect 1954 -9038 1971 -9011
rect 1888 -9038 1905 -9011
rect 1162 -9109 1179 -9082
rect 1096 -9109 1113 -9082
rect 1294 -9109 1311 -9082
rect 1228 -9109 1245 -9082
rect 1426 -9109 1443 -9082
rect 1360 -9109 1377 -9082
rect 1558 -9109 1575 -9082
rect 1492 -9109 1509 -9082
rect 1690 -9109 1707 -9082
rect 1624 -9109 1641 -9082
rect 1822 -9109 1839 -9082
rect 1756 -9109 1773 -9082
rect 1954 -9109 1971 -9082
rect 1954 -9109 1971 -9082
rect 1888 -9109 1905 -9082
rect 8 200 25 227
rect 64 200 81 227
rect 140 200 157 227
rect 196 200 213 227
rect 272 200 289 227
rect 328 200 345 227
rect 404 200 421 227
rect 460 200 477 227
rect 536 200 553 227
rect 592 200 609 227
rect 668 200 685 227
rect 724 200 741 227
rect 800 200 817 227
rect 856 200 873 227
rect 1129 200 1146 227
rect 1073 200 1090 227
rect 1261 200 1278 227
rect 1205 200 1222 227
rect 1393 200 1410 227
rect 1337 200 1354 227
rect 1525 200 1542 227
rect 1469 200 1486 227
rect 1657 200 1674 227
rect 1601 200 1618 227
rect 1789 200 1806 227
rect 1733 200 1750 227
rect 1921 200 1938 227
rect 1865 200 1882 227
<< nsubdiff >>
rect -89 27 1934 55
rect -91 -9133 -63 5
<< nsubdiffcont >>
rect -77 27 1922 55
rect -91 -9121 -63 -7
<< psubdiff >>
rect -89 262 1934 290
rect 1034 -9183 1967 -9155
<< psubdiffcont >>
rect -77 262 1922 290
rect 1046 -9183 1955 -9155
<< labels >>
flabel metal1 1946 -100 1979 -57 0 FreeSerif 160 0 0 0 word0
port 100 nsew
flabel metal1 1946 -171 1979 -128 0 FreeSerif 160 0 0 0 word1
port 101 nsew
flabel metal1 1946 -242 1979 -199 0 FreeSerif 160 0 0 0 word2
port 102 nsew
flabel metal1 1946 -313 1979 -270 0 FreeSerif 160 0 0 0 word3
port 103 nsew
flabel metal1 1946 -384 1979 -341 0 FreeSerif 160 0 0 0 word4
port 104 nsew
flabel metal1 1946 -455 1979 -412 0 FreeSerif 160 0 0 0 word5
port 105 nsew
flabel metal1 1946 -526 1979 -483 0 FreeSerif 160 0 0 0 word6
port 106 nsew
flabel metal1 1946 -597 1979 -554 0 FreeSerif 160 0 0 0 word7
port 107 nsew
flabel metal1 1946 -668 1979 -625 0 FreeSerif 160 0 0 0 word8
port 108 nsew
flabel metal1 1946 -739 1979 -696 0 FreeSerif 160 0 0 0 word9
port 109 nsew
flabel metal1 1946 -810 1979 -767 0 FreeSerif 160 0 0 0 word10
port 110 nsew
flabel metal1 1946 -881 1979 -838 0 FreeSerif 160 0 0 0 word11
port 111 nsew
flabel metal1 1946 -952 1979 -909 0 FreeSerif 160 0 0 0 word12
port 112 nsew
flabel metal1 1946 -1023 1979 -980 0 FreeSerif 160 0 0 0 word13
port 113 nsew
flabel metal1 1946 -1094 1979 -1051 0 FreeSerif 160 0 0 0 word14
port 114 nsew
flabel metal1 1946 -1165 1979 -1122 0 FreeSerif 160 0 0 0 word15
port 115 nsew
flabel metal1 1946 -1236 1979 -1193 0 FreeSerif 160 0 0 0 word16
port 116 nsew
flabel metal1 1946 -1307 1979 -1264 0 FreeSerif 160 0 0 0 word17
port 117 nsew
flabel metal1 1946 -1378 1979 -1335 0 FreeSerif 160 0 0 0 word18
port 118 nsew
flabel metal1 1946 -1449 1979 -1406 0 FreeSerif 160 0 0 0 word19
port 119 nsew
flabel metal1 1946 -1520 1979 -1477 0 FreeSerif 160 0 0 0 word20
port 120 nsew
flabel metal1 1946 -1591 1979 -1548 0 FreeSerif 160 0 0 0 word21
port 121 nsew
flabel metal1 1946 -1662 1979 -1619 0 FreeSerif 160 0 0 0 word22
port 122 nsew
flabel metal1 1946 -1733 1979 -1690 0 FreeSerif 160 0 0 0 word23
port 123 nsew
flabel metal1 1946 -1804 1979 -1761 0 FreeSerif 160 0 0 0 word24
port 124 nsew
flabel metal1 1946 -1875 1979 -1832 0 FreeSerif 160 0 0 0 word25
port 125 nsew
flabel metal1 1946 -1946 1979 -1903 0 FreeSerif 160 0 0 0 word26
port 126 nsew
flabel metal1 1946 -2017 1979 -1974 0 FreeSerif 160 0 0 0 word27
port 127 nsew
flabel metal1 1946 -2088 1979 -2045 0 FreeSerif 160 0 0 0 word28
port 128 nsew
flabel metal1 1946 -2159 1979 -2116 0 FreeSerif 160 0 0 0 word29
port 129 nsew
flabel metal1 1946 -2230 1979 -2187 0 FreeSerif 160 0 0 0 word30
port 130 nsew
flabel metal1 1946 -2301 1979 -2258 0 FreeSerif 160 0 0 0 word31
port 131 nsew
flabel metal1 1946 -2372 1979 -2329 0 FreeSerif 160 0 0 0 word32
port 132 nsew
flabel metal1 1946 -2443 1979 -2400 0 FreeSerif 160 0 0 0 word33
port 133 nsew
flabel metal1 1946 -2514 1979 -2471 0 FreeSerif 160 0 0 0 word34
port 134 nsew
flabel metal1 1946 -2585 1979 -2542 0 FreeSerif 160 0 0 0 word35
port 135 nsew
flabel metal1 1946 -2656 1979 -2613 0 FreeSerif 160 0 0 0 word36
port 136 nsew
flabel metal1 1946 -2727 1979 -2684 0 FreeSerif 160 0 0 0 word37
port 137 nsew
flabel metal1 1946 -2798 1979 -2755 0 FreeSerif 160 0 0 0 word38
port 138 nsew
flabel metal1 1946 -2869 1979 -2826 0 FreeSerif 160 0 0 0 word39
port 139 nsew
flabel metal1 1946 -2940 1979 -2897 0 FreeSerif 160 0 0 0 word40
port 140 nsew
flabel metal1 1946 -3011 1979 -2968 0 FreeSerif 160 0 0 0 word41
port 141 nsew
flabel metal1 1946 -3082 1979 -3039 0 FreeSerif 160 0 0 0 word42
port 142 nsew
flabel metal1 1946 -3153 1979 -3110 0 FreeSerif 160 0 0 0 word43
port 143 nsew
flabel metal1 1946 -3224 1979 -3181 0 FreeSerif 160 0 0 0 word44
port 144 nsew
flabel metal1 1946 -3295 1979 -3252 0 FreeSerif 160 0 0 0 word45
port 145 nsew
flabel metal1 1946 -3366 1979 -3323 0 FreeSerif 160 0 0 0 word46
port 146 nsew
flabel metal1 1946 -3437 1979 -3394 0 FreeSerif 160 0 0 0 word47
port 147 nsew
flabel metal1 1946 -3508 1979 -3465 0 FreeSerif 160 0 0 0 word48
port 148 nsew
flabel metal1 1946 -3579 1979 -3536 0 FreeSerif 160 0 0 0 word49
port 149 nsew
flabel metal1 1946 -3650 1979 -3607 0 FreeSerif 160 0 0 0 word50
port 150 nsew
flabel metal1 1946 -3721 1979 -3678 0 FreeSerif 160 0 0 0 word51
port 151 nsew
flabel metal1 1946 -3792 1979 -3749 0 FreeSerif 160 0 0 0 word52
port 152 nsew
flabel metal1 1946 -3863 1979 -3820 0 FreeSerif 160 0 0 0 word53
port 153 nsew
flabel metal1 1946 -3934 1979 -3891 0 FreeSerif 160 0 0 0 word54
port 154 nsew
flabel metal1 1946 -4005 1979 -3962 0 FreeSerif 160 0 0 0 word55
port 155 nsew
flabel metal1 1946 -4076 1979 -4033 0 FreeSerif 160 0 0 0 word56
port 156 nsew
flabel metal1 1946 -4147 1979 -4104 0 FreeSerif 160 0 0 0 word57
port 157 nsew
flabel metal1 1946 -4218 1979 -4175 0 FreeSerif 160 0 0 0 word58
port 158 nsew
flabel metal1 1946 -4289 1979 -4246 0 FreeSerif 160 0 0 0 word59
port 159 nsew
flabel metal1 1946 -4360 1979 -4317 0 FreeSerif 160 0 0 0 word60
port 160 nsew
flabel metal1 1946 -4431 1979 -4388 0 FreeSerif 160 0 0 0 word61
port 161 nsew
flabel metal1 1946 -4502 1979 -4459 0 FreeSerif 160 0 0 0 word62
port 162 nsew
flabel metal1 1946 -4573 1979 -4530 0 FreeSerif 160 0 0 0 word63
port 163 nsew
flabel metal1 1946 -4644 1979 -4601 0 FreeSerif 160 0 0 0 word64
port 164 nsew
flabel metal1 1946 -4715 1979 -4672 0 FreeSerif 160 0 0 0 word65
port 165 nsew
flabel metal1 1946 -4786 1979 -4743 0 FreeSerif 160 0 0 0 word66
port 166 nsew
flabel metal1 1946 -4857 1979 -4814 0 FreeSerif 160 0 0 0 word67
port 167 nsew
flabel metal1 1946 -4928 1979 -4885 0 FreeSerif 160 0 0 0 word68
port 168 nsew
flabel metal1 1946 -4999 1979 -4956 0 FreeSerif 160 0 0 0 word69
port 169 nsew
flabel metal1 1946 -5070 1979 -5027 0 FreeSerif 160 0 0 0 word70
port 170 nsew
flabel metal1 1946 -5141 1979 -5098 0 FreeSerif 160 0 0 0 word71
port 171 nsew
flabel metal1 1946 -5212 1979 -5169 0 FreeSerif 160 0 0 0 word72
port 172 nsew
flabel metal1 1946 -5283 1979 -5240 0 FreeSerif 160 0 0 0 word73
port 173 nsew
flabel metal1 1946 -5354 1979 -5311 0 FreeSerif 160 0 0 0 word74
port 174 nsew
flabel metal1 1946 -5425 1979 -5382 0 FreeSerif 160 0 0 0 word75
port 175 nsew
flabel metal1 1946 -5496 1979 -5453 0 FreeSerif 160 0 0 0 word76
port 176 nsew
flabel metal1 1946 -5567 1979 -5524 0 FreeSerif 160 0 0 0 word77
port 177 nsew
flabel metal1 1946 -5638 1979 -5595 0 FreeSerif 160 0 0 0 word78
port 178 nsew
flabel metal1 1946 -5709 1979 -5666 0 FreeSerif 160 0 0 0 word79
port 179 nsew
flabel metal1 1946 -5780 1979 -5737 0 FreeSerif 160 0 0 0 word80
port 180 nsew
flabel metal1 1946 -5851 1979 -5808 0 FreeSerif 160 0 0 0 word81
port 181 nsew
flabel metal1 1946 -5922 1979 -5879 0 FreeSerif 160 0 0 0 word82
port 182 nsew
flabel metal1 1946 -5993 1979 -5950 0 FreeSerif 160 0 0 0 word83
port 183 nsew
flabel metal1 1946 -6064 1979 -6021 0 FreeSerif 160 0 0 0 word84
port 184 nsew
flabel metal1 1946 -6135 1979 -6092 0 FreeSerif 160 0 0 0 word85
port 185 nsew
flabel metal1 1946 -6206 1979 -6163 0 FreeSerif 160 0 0 0 word86
port 186 nsew
flabel metal1 1946 -6277 1979 -6234 0 FreeSerif 160 0 0 0 word87
port 187 nsew
flabel metal1 1946 -6348 1979 -6305 0 FreeSerif 160 0 0 0 word88
port 188 nsew
flabel metal1 1946 -6419 1979 -6376 0 FreeSerif 160 0 0 0 word89
port 189 nsew
flabel metal1 1946 -6490 1979 -6447 0 FreeSerif 160 0 0 0 word90
port 190 nsew
flabel metal1 1946 -6561 1979 -6518 0 FreeSerif 160 0 0 0 word91
port 191 nsew
flabel metal1 1946 -6632 1979 -6589 0 FreeSerif 160 0 0 0 word92
port 192 nsew
flabel metal1 1946 -6703 1979 -6660 0 FreeSerif 160 0 0 0 word93
port 193 nsew
flabel metal1 1946 -6774 1979 -6731 0 FreeSerif 160 0 0 0 word94
port 194 nsew
flabel metal1 1946 -6845 1979 -6802 0 FreeSerif 160 0 0 0 word95
port 195 nsew
flabel metal1 1946 -6916 1979 -6873 0 FreeSerif 160 0 0 0 word96
port 196 nsew
flabel metal1 1946 -6987 1979 -6944 0 FreeSerif 160 0 0 0 word97
port 197 nsew
flabel metal1 1946 -7058 1979 -7015 0 FreeSerif 160 0 0 0 word98
port 198 nsew
flabel metal1 1946 -7129 1979 -7086 0 FreeSerif 160 0 0 0 word99
port 199 nsew
flabel metal1 1946 -7200 1979 -7157 0 FreeSerif 160 0 0 0 word100
port 200 nsew
flabel metal1 1946 -7271 1979 -7228 0 FreeSerif 160 0 0 0 word101
port 201 nsew
flabel metal1 1946 -7342 1979 -7299 0 FreeSerif 160 0 0 0 word102
port 202 nsew
flabel metal1 1946 -7413 1979 -7370 0 FreeSerif 160 0 0 0 word103
port 203 nsew
flabel metal1 1946 -7484 1979 -7441 0 FreeSerif 160 0 0 0 word104
port 204 nsew
flabel metal1 1946 -7555 1979 -7512 0 FreeSerif 160 0 0 0 word105
port 205 nsew
flabel metal1 1946 -7626 1979 -7583 0 FreeSerif 160 0 0 0 word106
port 206 nsew
flabel metal1 1946 -7697 1979 -7654 0 FreeSerif 160 0 0 0 word107
port 207 nsew
flabel metal1 1946 -7768 1979 -7725 0 FreeSerif 160 0 0 0 word108
port 208 nsew
flabel metal1 1946 -7839 1979 -7796 0 FreeSerif 160 0 0 0 word109
port 209 nsew
flabel metal1 1946 -7910 1979 -7867 0 FreeSerif 160 0 0 0 word110
port 210 nsew
flabel metal1 1946 -7981 1979 -7938 0 FreeSerif 160 0 0 0 word111
port 211 nsew
flabel metal1 1946 -8052 1979 -8009 0 FreeSerif 160 0 0 0 word112
port 212 nsew
flabel metal1 1946 -8123 1979 -8080 0 FreeSerif 160 0 0 0 word113
port 213 nsew
flabel metal1 1946 -8194 1979 -8151 0 FreeSerif 160 0 0 0 word114
port 214 nsew
flabel metal1 1946 -8265 1979 -8222 0 FreeSerif 160 0 0 0 word115
port 215 nsew
flabel metal1 1946 -8336 1979 -8293 0 FreeSerif 160 0 0 0 word116
port 216 nsew
flabel metal1 1946 -8407 1979 -8364 0 FreeSerif 160 0 0 0 word117
port 217 nsew
flabel metal1 1946 -8478 1979 -8435 0 FreeSerif 160 0 0 0 word118
port 218 nsew
flabel metal1 1946 -8549 1979 -8506 0 FreeSerif 160 0 0 0 word119
port 219 nsew
flabel metal1 1946 -8620 1979 -8577 0 FreeSerif 160 0 0 0 word120
port 220 nsew
flabel metal1 1946 -8691 1979 -8648 0 FreeSerif 160 0 0 0 word121
port 221 nsew
flabel metal1 1946 -8762 1979 -8719 0 FreeSerif 160 0 0 0 word122
port 222 nsew
flabel metal1 1946 -8833 1979 -8790 0 FreeSerif 160 0 0 0 word123
port 223 nsew
flabel metal1 1946 -8904 1979 -8861 0 FreeSerif 160 0 0 0 word124
port 224 nsew
flabel metal1 1946 -8975 1979 -8932 0 FreeSerif 160 0 0 0 word125
port 225 nsew
flabel metal1 1946 -9046 1979 -9003 0 FreeSerif 160 0 0 0 word126
port 226 nsew
flabel metal1 1946 -9117 1979 -9074 0 FreeSerif 160 0 0 0 word127
port 227 nsew
flabel locali -101 -9145 -53 17 0 FreeSerif 160 0 0 0 VDD!
port 228 nsew
flabel locali 2019 -9145 2059 300 0 FreeSerif 160 0 0 0 GND!
port 229 nsew
flabel metal2 891 142 924 175 0 FreeSerif 160 0 0 0 A0
port 19 nsew
flabel metal2 759 189 792 222 0 FreeSerif 160 0 0 0 A1
port 20 nsew
flabel metal2 627 236 660 269 0 FreeSerif 160 0 0 0 A2
port 21 nsew
flabel metal2 495 283 528 316 0 FreeSerif 160 0 0 0 A3
port 22 nsew
flabel metal2 363 330 396 363 0 FreeSerif 160 0 0 0 A4
port 23 nsew
flabel metal2 231 377 264 410 0 FreeSerif 160 0 0 0 A5
port 24 nsew
flabel metal2 99 424 132 457 0 FreeSerif 160 0 0 0 A6
port 25 nsew
<< end >>