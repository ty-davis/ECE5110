magic
tech sky130A
timestamp 1741799890
<< nwell >>
rect 3 197 189 488
<< nmos >>
rect 72 65 87 115
rect 108 65 123 115
<< pmos >>
rect 72 315 87 415
rect 108 315 123 415
<< ndiff >>
rect 36 107 72 115
rect 36 73 44 107
rect 61 73 72 107
rect 36 65 72 73
rect 87 65 108 115
rect 123 107 159 115
rect 123 73 134 107
rect 151 73 159 107
rect 123 65 159 73
<< pdiff >>
rect 36 407 72 415
rect 36 323 44 407
rect 61 323 72 407
rect 36 315 72 323
rect 87 315 108 415
rect 123 407 159 415
rect 123 323 134 407
rect 151 323 159 407
rect 123 315 159 323
<< ndiffc >>
rect 44 73 61 107
rect 134 73 151 107
<< pdiffc >>
rect 44 323 61 407
rect 134 323 151 407
<< psubdiff >>
rect 5 10 17 38
rect 175 10 187 38
<< nsubdiff >>
rect 21 442 33 470
rect 159 442 171 470
<< psubdiffcont >>
rect 17 10 175 38
<< nsubdiffcont >>
rect 33 442 159 470
<< poly >>
rect 72 415 87 428
rect 108 415 123 428
rect 72 298 87 315
rect 33 290 87 298
rect 33 273 41 290
rect 58 283 87 290
rect 58 273 66 283
rect 33 265 66 273
rect 36 138 52 265
rect 108 246 123 315
rect 75 238 123 246
rect 75 221 83 238
rect 100 231 123 238
rect 100 221 108 231
rect 75 213 108 221
rect 75 184 108 192
rect 75 167 83 184
rect 100 167 123 184
rect 75 159 123 167
rect 36 123 87 138
rect 72 115 87 123
rect 108 115 123 159
rect 72 52 87 65
rect 108 52 123 65
<< polycont >>
rect 41 273 58 290
rect 83 221 100 238
rect 83 167 100 184
<< locali >>
rect 5 470 187 480
rect 5 442 33 470
rect 159 442 187 470
rect 5 432 187 442
rect 36 407 69 432
rect 36 323 44 407
rect 61 323 69 407
rect 36 315 69 323
rect 126 407 159 415
rect 126 323 134 407
rect 151 323 159 407
rect 33 290 66 298
rect 33 273 41 290
rect 58 273 66 290
rect 33 265 66 273
rect 75 238 108 246
rect 75 221 83 238
rect 100 221 108 238
rect 75 213 108 221
rect 75 184 108 192
rect 75 167 83 184
rect 100 167 108 184
rect 75 159 108 167
rect 36 107 69 115
rect 36 73 44 107
rect 61 73 69 107
rect 36 48 69 73
rect 126 107 159 323
rect 126 73 134 107
rect 151 73 159 107
rect 126 65 159 73
rect 5 38 187 48
rect 5 10 17 38
rect 175 10 187 38
rect 5 0 187 10
<< labels >>
flabel ndiff 72 90 72 90 1 FreeSerif 8 0 0 0 S$
flabel pdiff 72 365 72 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 108 365 108 365 1 FreeSerif 8 0 0 0 S$
flabel ndiff 108 90 108 90 1 FreeSerif 8 0 0 0 S$
flabel locali 126 115 159 315 0 FreeSerif 80 0 0 0 Y
port 5 nsew
flabel locali 75 159 108 192 0 FreeSerif 80 0 0 0 EN
port 8 nsew
flabel locali 75 213 108 246 0 FreeSerif 80 0 0 0 ~EN
port 9 nsew
flabel locali 33 265 66 298 0 FreeSerif 80 0 0 0 A
port 4 nsew
flabel locali 5 432 187 480 0 FreeSerif 80 0 0 0 VDD!
port 2 nsew
flabel locali 5 0 187 48 0 FreeSerif 80 0 0 0 GND!
port 3 nsew
<< end >>
