magic
tech sky130A
magscale 1 2
timestamp 1745497054
<< error_s >>
rect 60 145672 166 145682
<< nwell >>
rect -816 119516 -782 119552
rect 0 80 2914 118
<< locali >>
rect -114 146128 84 146176
rect -974 145854 -926 145860
rect -974 145818 -968 145854
rect -932 145818 -926 145854
rect -974 145626 -926 145818
rect -114 145628 -66 146128
rect 5758 146042 5814 146048
rect 5758 145998 5764 146042
rect 5808 145998 5814 146042
rect 36 145700 84 145818
rect 5758 145732 5814 145998
rect 6028 145992 6114 146048
rect 5660 145676 5814 145732
rect 5860 145626 6040 145706
rect -577 119909 -511 120090
rect -830 119563 -770 119564
rect -619 119563 -553 119782
rect -839 119552 -553 119563
rect -839 119516 -820 119552
rect -782 119516 -553 119552
rect -839 119504 -553 119516
rect 50 -84 106 140
rect 50 -128 56 -84
rect 100 -128 106 -84
rect 50 -134 106 -128
rect 5270 -924 5366 18
rect 5598 -134 5704 -78
rect 5828 -674 5894 -472
rect 6136 -674 6202 -472
rect 6444 -674 6510 -472
rect 6752 -564 6818 -362
rect 7060 -584 7126 -382
rect 7368 -592 7434 -390
rect 7676 -594 7742 -392
rect 7984 -598 8050 -396
rect 5270 -1020 5670 -924
<< viali >>
rect -968 145818 -932 145854
rect 5764 145998 5808 146042
rect 36 145818 84 145854
rect 5984 145992 6028 146048
rect 6015 145436 6032 145486
rect 6015 145294 6032 145344
rect 6015 145152 6032 145202
rect 6015 145010 6032 145060
rect 6015 144868 6032 144918
rect 6015 144726 6032 144776
rect 6015 144584 6032 144634
rect 6015 144442 6032 144492
rect 6015 144300 6032 144350
rect 6015 144158 6032 144208
rect 6015 144016 6032 144066
rect 6015 143874 6032 143924
rect 6015 143732 6032 143782
rect 6015 143590 6032 143640
rect 6015 143448 6032 143498
rect 6015 143306 6032 143356
rect 6015 143164 6032 143214
rect 6015 143022 6032 143072
rect 6015 142880 6032 142930
rect 6015 142738 6032 142788
rect 6015 142596 6032 142646
rect 6015 142454 6032 142504
rect 6015 142312 6032 142362
rect 6015 142170 6032 142220
rect 6015 142028 6032 142078
rect 6015 141886 6032 141936
rect 6015 141744 6032 141794
rect 6015 141602 6032 141652
rect 6015 141460 6032 141510
rect 6015 141318 6032 141368
rect 6015 141176 6032 141226
rect 6015 141034 6032 141084
rect 6015 140892 6032 140942
rect 6015 140750 6032 140800
rect 6015 140608 6032 140658
rect 6015 140466 6032 140516
rect 6015 140324 6032 140374
rect 6015 140182 6032 140232
rect 6015 140040 6032 140090
rect 6015 139898 6032 139948
rect 6015 139756 6032 139806
rect 6015 139614 6032 139664
rect 6015 139472 6032 139522
rect 6015 139330 6032 139380
rect 6015 139188 6032 139238
rect 6015 139046 6032 139096
rect 6015 138904 6032 138954
rect 6015 138762 6032 138812
rect 6015 138620 6032 138670
rect 6015 138478 6032 138528
rect 6015 138336 6032 138386
rect 6015 138194 6032 138244
rect 6015 138052 6032 138102
rect 6015 137910 6032 137960
rect 6015 137768 6032 137818
rect 6015 137626 6032 137676
rect 6015 137484 6032 137534
rect 6015 137342 6032 137392
rect 6015 137200 6032 137250
rect 6015 137058 6032 137108
rect 6015 136916 6032 136966
rect 6015 136774 6032 136824
rect 6015 136632 6032 136682
rect 6015 136490 6032 136540
rect 6015 136348 6032 136398
rect 6015 136206 6032 136256
rect 6015 136064 6032 136114
rect 6015 135922 6032 135972
rect 6015 135780 6032 135830
rect 6015 135638 6032 135688
rect 6015 135496 6032 135546
rect 6015 135354 6032 135404
rect 6015 135212 6032 135262
rect 6015 135070 6032 135120
rect 6015 134928 6032 134978
rect 6015 134786 6032 134836
rect 6015 134644 6032 134694
rect 6015 134502 6032 134552
rect 6015 134360 6032 134410
rect 6015 134218 6032 134268
rect 6015 134076 6032 134126
rect 6015 133934 6032 133984
rect 6015 133792 6032 133842
rect 6015 133650 6032 133700
rect 6015 133508 6032 133558
rect 6015 133366 6032 133416
rect 6015 133224 6032 133274
rect 6015 133082 6032 133132
rect 6015 132940 6032 132990
rect 6015 132798 6032 132848
rect 6015 132656 6032 132706
rect 6015 132514 6032 132564
rect 6015 132372 6032 132422
rect 6015 132230 6032 132280
rect 6015 132088 6032 132138
rect 6015 131946 6032 131996
rect 6015 131804 6032 131854
rect 6015 131662 6032 131712
rect 6015 131520 6032 131570
rect 6015 131378 6032 131428
rect 6015 131236 6032 131286
rect 6015 131094 6032 131144
rect 6015 130952 6032 131002
rect 6015 130810 6032 130860
rect 6015 130668 6032 130718
rect 6015 130526 6032 130576
rect 6015 130384 6032 130434
rect 6015 130242 6032 130292
rect 6015 130100 6032 130150
rect 6015 129958 6032 130008
rect 6015 129816 6032 129866
rect 6015 129674 6032 129724
rect 6015 129532 6032 129582
rect 6015 129390 6032 129440
rect 6015 129248 6032 129298
rect 6015 129106 6032 129156
rect 6015 128964 6032 129014
rect 6015 128822 6032 128872
rect 6015 128680 6032 128730
rect 6015 128538 6032 128588
rect 6015 128396 6032 128446
rect 6015 128254 6032 128304
rect 6015 128112 6032 128162
rect 6015 127970 6032 128020
rect 6015 127828 6032 127878
rect 6015 127686 6032 127736
rect 6015 127544 6032 127594
rect 6015 127402 6032 127452
rect 6015 127260 6032 127310
rect 6015 127118 6032 127168
rect 6015 126976 6032 127026
rect 6015 126834 6032 126884
rect 6015 126692 6032 126742
rect 6015 126550 6032 126600
rect 6015 126408 6032 126458
rect 6015 126266 6032 126316
rect 6015 126124 6032 126174
rect 6015 125982 6032 126032
rect 6015 125840 6032 125890
rect 6015 125698 6032 125748
rect 6015 125556 6032 125606
rect 6015 125414 6032 125464
rect 6015 125272 6032 125322
rect 6015 125130 6032 125180
rect 6015 124988 6032 125038
rect 6015 124846 6032 124896
rect 6015 124704 6032 124754
rect 6015 124562 6032 124612
rect 6015 124420 6032 124470
rect 6015 124278 6032 124328
rect 6015 124136 6032 124186
rect 6015 123994 6032 124044
rect 6015 123852 6032 123902
rect 6015 123710 6032 123760
rect 6015 123568 6032 123618
rect 6015 123426 6032 123476
rect 6015 123284 6032 123334
rect 6015 123142 6032 123192
rect 6015 123000 6032 123050
rect 6015 122858 6032 122908
rect 6015 122716 6032 122766
rect 6015 122574 6032 122624
rect 6015 122432 6032 122482
rect 6015 122290 6032 122340
rect 6015 122148 6032 122198
rect 6015 122006 6032 122056
rect 6015 121864 6032 121914
rect 6015 121722 6032 121772
rect 6015 121580 6032 121630
rect 6015 121438 6032 121488
rect 6015 121296 6032 121346
rect 6015 121154 6032 121204
rect 6015 121012 6032 121062
rect 6015 120870 6032 120920
rect 6015 120728 6032 120778
rect 6015 120586 6032 120636
rect 6015 120444 6032 120494
rect 6015 120302 6032 120352
rect 6015 120160 6032 120210
rect 6015 120018 6032 120068
rect -390 119936 -348 119976
rect -577 119855 -511 119909
rect 6015 119876 6032 119926
rect 6015 119734 6032 119784
rect -388 119628 -352 119670
rect 6015 119592 6032 119642
rect -820 119516 -782 119552
rect -518 119462 -452 119528
rect 6015 119450 6032 119500
rect 6015 119308 6032 119358
rect -533 119223 -479 119277
rect -533 119115 -479 119169
rect 6015 119166 6032 119216
rect 6015 119024 6032 119074
rect 6015 118882 6032 118932
rect -631 118767 -577 118821
rect 6015 118740 6032 118790
rect 6015 118598 6032 118648
rect 6015 118456 6032 118506
rect -613 118365 -559 118419
rect 6015 118314 6032 118364
rect -631 118131 -577 118185
rect 6015 118172 6032 118222
rect 6015 118030 6032 118080
rect 6015 117888 6032 117938
rect -621 117735 -551 117805
rect 6015 117746 6032 117796
rect 6015 117604 6032 117654
rect 6015 117462 6032 117512
rect -471 117316 -417 117370
rect 6015 117320 6032 117370
rect 6015 117178 6032 117228
rect 6015 117036 6032 117086
rect 6015 116894 6032 116944
rect 6015 116752 6032 116802
rect 6015 116610 6032 116660
rect 6015 116468 6032 116518
rect 6015 116326 6032 116376
rect 6015 116184 6032 116234
rect 6015 116042 6032 116092
rect 6015 115900 6032 115950
rect 6015 115758 6032 115808
rect 6015 115616 6032 115666
rect 6015 115474 6032 115524
rect 6015 115332 6032 115382
rect 6015 115190 6032 115240
rect 6015 115048 6032 115098
rect 6015 114906 6032 114956
rect 6015 114764 6032 114814
rect 6015 114622 6032 114672
rect 6015 114480 6032 114530
rect 6015 114338 6032 114388
rect 6015 114196 6032 114246
rect 6015 114054 6032 114104
rect 6015 113912 6032 113962
rect 6015 113770 6032 113820
rect 6015 113628 6032 113678
rect 6015 113486 6032 113536
rect 6015 113344 6032 113394
rect 6015 113202 6032 113252
rect 6015 113060 6032 113110
rect 6015 112918 6032 112968
rect 6015 112776 6032 112826
rect 6015 112634 6032 112684
rect 6015 112492 6032 112542
rect 6015 112350 6032 112400
rect 6015 112208 6032 112258
rect 6015 112066 6032 112116
rect 6015 111924 6032 111974
rect 6015 111782 6032 111832
rect 6015 111640 6032 111690
rect 6015 111498 6032 111548
rect 6015 111356 6032 111406
rect 6015 111214 6032 111264
rect 6015 111072 6032 111122
rect 6015 110930 6032 110980
rect 6015 110788 6032 110838
rect 6015 110646 6032 110696
rect 6015 110504 6032 110554
rect 6015 110362 6032 110412
rect 6015 110220 6032 110270
rect 6015 110078 6032 110128
rect 6015 109936 6032 109986
rect 6015 109794 6032 109844
rect 6015 109652 6032 109702
rect 6015 109510 6032 109560
rect 6015 109368 6032 109418
rect 6015 109226 6032 109276
rect 6015 109084 6032 109134
rect 6015 108942 6032 108992
rect 6015 108800 6032 108850
rect 6015 108658 6032 108708
rect 6015 108516 6032 108566
rect 6015 108374 6032 108424
rect 6015 108232 6032 108282
rect 6015 108090 6032 108140
rect 6015 107948 6032 107998
rect 6015 107806 6032 107856
rect 6015 107664 6032 107714
rect 6015 107522 6032 107572
rect 6015 107380 6032 107430
rect 6015 107238 6032 107288
rect 6015 107096 6032 107146
rect 6015 106954 6032 107004
rect 6015 106812 6032 106862
rect 6015 106670 6032 106720
rect 6015 106528 6032 106578
rect 6015 106386 6032 106436
rect 6015 106244 6032 106294
rect 6015 106102 6032 106152
rect 6015 105960 6032 106010
rect 6015 105818 6032 105868
rect 6015 105676 6032 105726
rect 6015 105534 6032 105584
rect 6015 105392 6032 105442
rect 6015 105250 6032 105300
rect 6015 105108 6032 105158
rect 6015 104966 6032 105016
rect 6015 104824 6032 104874
rect 6015 104682 6032 104732
rect 6015 104540 6032 104590
rect 6015 104398 6032 104448
rect 6015 104256 6032 104306
rect 6015 104114 6032 104164
rect 6015 103972 6032 104022
rect 6015 103830 6032 103880
rect 6015 103688 6032 103738
rect 6015 103546 6032 103596
rect 6015 103404 6032 103454
rect 6015 103262 6032 103312
rect 6015 103120 6032 103170
rect 6015 102978 6032 103028
rect 6015 102836 6032 102886
rect 6015 102694 6032 102744
rect 6015 102552 6032 102602
rect 6015 102410 6032 102460
rect 6015 102268 6032 102318
rect 6015 102126 6032 102176
rect 6015 101984 6032 102034
rect 6015 101842 6032 101892
rect 6015 101700 6032 101750
rect 6015 101558 6032 101608
rect 6015 101416 6032 101466
rect 6015 101274 6032 101324
rect 6015 101132 6032 101182
rect 6015 100990 6032 101040
rect 6015 100848 6032 100898
rect 6015 100706 6032 100756
rect 6015 100564 6032 100614
rect 6015 100422 6032 100472
rect 6015 100280 6032 100330
rect 6015 100138 6032 100188
rect 6015 99996 6032 100046
rect 6015 99854 6032 99904
rect 6015 99712 6032 99762
rect 6015 99570 6032 99620
rect 6015 99428 6032 99478
rect 6015 99286 6032 99336
rect 6015 99144 6032 99194
rect 6015 99002 6032 99052
rect 6015 98860 6032 98910
rect 6015 98718 6032 98768
rect 6015 98576 6032 98626
rect 6015 98434 6032 98484
rect 6015 98292 6032 98342
rect 6015 98150 6032 98200
rect 6015 98008 6032 98058
rect 6015 97866 6032 97916
rect 6015 97724 6032 97774
rect 6015 97582 6032 97632
rect 6015 97440 6032 97490
rect 6015 97298 6032 97348
rect 6015 97156 6032 97206
rect 6015 97014 6032 97064
rect 6015 96872 6032 96922
rect 6015 96730 6032 96780
rect 6015 96588 6032 96638
rect 6015 96446 6032 96496
rect 6015 96304 6032 96354
rect 6015 96162 6032 96212
rect 6015 96020 6032 96070
rect 6015 95878 6032 95928
rect 6015 95736 6032 95786
rect 6015 95594 6032 95644
rect 6015 95452 6032 95502
rect 6015 95310 6032 95360
rect 6015 95168 6032 95218
rect 6015 95026 6032 95076
rect 6015 94884 6032 94934
rect 6015 94742 6032 94792
rect 6015 94600 6032 94650
rect 6015 94458 6032 94508
rect 6015 94316 6032 94366
rect 6015 94174 6032 94224
rect 6015 94032 6032 94082
rect 6015 93890 6032 93940
rect 6015 93748 6032 93798
rect 6015 93606 6032 93656
rect 6015 93464 6032 93514
rect 6015 93322 6032 93372
rect 6015 93180 6032 93230
rect 6015 93038 6032 93088
rect 6015 92896 6032 92946
rect 6015 92754 6032 92804
rect 6015 92612 6032 92662
rect 6015 92470 6032 92520
rect 6015 92328 6032 92378
rect 6015 92186 6032 92236
rect 6015 92044 6032 92094
rect 6015 91902 6032 91952
rect 6015 91760 6032 91810
rect 6015 91618 6032 91668
rect 6015 91476 6032 91526
rect 6015 91334 6032 91384
rect 6015 91192 6032 91242
rect 6015 91050 6032 91100
rect 6015 90908 6032 90958
rect 6015 90766 6032 90816
rect 6015 90624 6032 90674
rect 6015 90482 6032 90532
rect 6015 90340 6032 90390
rect 6015 90198 6032 90248
rect 6015 90056 6032 90106
rect 6015 89914 6032 89964
rect 6015 89772 6032 89822
rect 6015 89630 6032 89680
rect 6015 89488 6032 89538
rect 6015 89346 6032 89396
rect 6015 89204 6032 89254
rect 6015 89062 6032 89112
rect 6015 88920 6032 88970
rect 6015 88778 6032 88828
rect 6015 88636 6032 88686
rect 6015 88494 6032 88544
rect 6015 88352 6032 88402
rect 6015 88210 6032 88260
rect 6015 88068 6032 88118
rect 6015 87926 6032 87976
rect 6015 87784 6032 87834
rect 6015 87642 6032 87692
rect 6015 87500 6032 87550
rect 6015 87358 6032 87408
rect 6015 87216 6032 87266
rect 6015 87074 6032 87124
rect 6015 86932 6032 86982
rect 6015 86790 6032 86840
rect 6015 86648 6032 86698
rect 6015 86506 6032 86556
rect 6015 86364 6032 86414
rect 6015 86222 6032 86272
rect 6015 86080 6032 86130
rect 6015 85938 6032 85988
rect 6015 85796 6032 85846
rect 6015 85654 6032 85704
rect 6015 85512 6032 85562
rect 6015 85370 6032 85420
rect 6015 85228 6032 85278
rect 6015 85086 6032 85136
rect 6015 84944 6032 84994
rect 6015 84802 6032 84852
rect 6015 84660 6032 84710
rect 6015 84518 6032 84568
rect 6015 84376 6032 84426
rect 6015 84234 6032 84284
rect 6015 84092 6032 84142
rect 6015 83950 6032 84000
rect 6015 83808 6032 83858
rect 6015 83666 6032 83716
rect 6015 83524 6032 83574
rect 6015 83382 6032 83432
rect 6015 83240 6032 83290
rect 6015 83098 6032 83148
rect 6015 82956 6032 83006
rect 6015 82814 6032 82864
rect 6015 82672 6032 82722
rect 6015 82530 6032 82580
rect 6015 82388 6032 82438
rect 6015 82246 6032 82296
rect 6015 82104 6032 82154
rect 6015 81962 6032 82012
rect 6015 81820 6032 81870
rect 6015 81678 6032 81728
rect 6015 81536 6032 81586
rect 6015 81394 6032 81444
rect 6015 81252 6032 81302
rect 6015 81110 6032 81160
rect 6015 80968 6032 81018
rect 6015 80826 6032 80876
rect 6015 80684 6032 80734
rect 6015 80542 6032 80592
rect 6015 80400 6032 80450
rect 6015 80258 6032 80308
rect 6015 80116 6032 80166
rect 6015 79974 6032 80024
rect 6015 79832 6032 79882
rect 6015 79690 6032 79740
rect 6015 79548 6032 79598
rect 6015 79406 6032 79456
rect 6015 79264 6032 79314
rect 6015 79122 6032 79172
rect 6015 78980 6032 79030
rect 6015 78838 6032 78888
rect 6015 78696 6032 78746
rect 6015 78554 6032 78604
rect 6015 78412 6032 78462
rect 6015 78270 6032 78320
rect 6015 78128 6032 78178
rect 6015 77986 6032 78036
rect 6015 77844 6032 77894
rect 6015 77702 6032 77752
rect 6015 77560 6032 77610
rect 6015 77418 6032 77468
rect 6015 77276 6032 77326
rect 6015 77134 6032 77184
rect 6015 76992 6032 77042
rect 6015 76850 6032 76900
rect 6015 76708 6032 76758
rect 6015 76566 6032 76616
rect 6015 76424 6032 76474
rect 6015 76282 6032 76332
rect 6015 76140 6032 76190
rect 6015 75998 6032 76048
rect 6015 75856 6032 75906
rect 6015 75714 6032 75764
rect 6015 75572 6032 75622
rect 6015 75430 6032 75480
rect 6015 75288 6032 75338
rect 6015 75146 6032 75196
rect 6015 75004 6032 75054
rect 6015 74862 6032 74912
rect 6015 74720 6032 74770
rect 6015 74578 6032 74628
rect 6015 74436 6032 74486
rect 6015 74294 6032 74344
rect 6015 74152 6032 74202
rect 6015 74010 6032 74060
rect 6015 73868 6032 73918
rect 6015 73726 6032 73776
rect 6015 73584 6032 73634
rect 6015 73442 6032 73492
rect 6015 73300 6032 73350
rect 6015 73158 6032 73208
rect 6015 73016 6032 73066
rect 6015 72874 6032 72924
rect 6015 72732 6032 72782
rect 6015 72590 6032 72640
rect 6015 72448 6032 72498
rect 6015 72306 6032 72356
rect 6015 72164 6032 72214
rect 6015 72022 6032 72072
rect 6015 71880 6032 71930
rect 6015 71738 6032 71788
rect 6015 71596 6032 71646
rect 6015 71454 6032 71504
rect 6015 71312 6032 71362
rect 6015 71170 6032 71220
rect 6015 71028 6032 71078
rect 6015 70886 6032 70936
rect 6015 70744 6032 70794
rect 6015 70602 6032 70652
rect 6015 70460 6032 70510
rect 6015 70318 6032 70368
rect 6015 70176 6032 70226
rect 6015 70034 6032 70084
rect 6015 69892 6032 69942
rect 6015 69750 6032 69800
rect 6015 69608 6032 69658
rect 6015 69466 6032 69516
rect 6015 69324 6032 69374
rect 6015 69182 6032 69232
rect 6015 69040 6032 69090
rect 6015 68898 6032 68948
rect 6015 68756 6032 68806
rect 6015 68614 6032 68664
rect 6015 68472 6032 68522
rect 6015 68330 6032 68380
rect 6015 68188 6032 68238
rect 6015 68046 6032 68096
rect 6015 67904 6032 67954
rect 6015 67762 6032 67812
rect 6015 67620 6032 67670
rect 6015 67478 6032 67528
rect 6015 67336 6032 67386
rect 6015 67194 6032 67244
rect 6015 67052 6032 67102
rect 6015 66910 6032 66960
rect 6015 66768 6032 66818
rect 6015 66626 6032 66676
rect 6015 66484 6032 66534
rect 6015 66342 6032 66392
rect 6015 66200 6032 66250
rect 6015 66058 6032 66108
rect 6015 65916 6032 65966
rect 6015 65774 6032 65824
rect 6015 65632 6032 65682
rect 6015 65490 6032 65540
rect 6015 65348 6032 65398
rect 6015 65206 6032 65256
rect 6015 65064 6032 65114
rect 6015 64922 6032 64972
rect 6015 64780 6032 64830
rect 6015 64638 6032 64688
rect 6015 64496 6032 64546
rect 6015 64354 6032 64404
rect 6015 64212 6032 64262
rect 6015 64070 6032 64120
rect 6015 63928 6032 63978
rect 6015 63786 6032 63836
rect 6015 63644 6032 63694
rect 6015 63502 6032 63552
rect 6015 63360 6032 63410
rect 6015 63218 6032 63268
rect 6015 63076 6032 63126
rect 6015 62934 6032 62984
rect 6015 62792 6032 62842
rect 6015 62650 6032 62700
rect 6015 62508 6032 62558
rect 6015 62366 6032 62416
rect 6015 62224 6032 62274
rect 6015 62082 6032 62132
rect 6015 61940 6032 61990
rect 6015 61798 6032 61848
rect 6015 61656 6032 61706
rect 6015 61514 6032 61564
rect 6015 61372 6032 61422
rect 6015 61230 6032 61280
rect 6015 61088 6032 61138
rect 6015 60946 6032 60996
rect 6015 60804 6032 60854
rect 6015 60662 6032 60712
rect 6015 60520 6032 60570
rect 6015 60378 6032 60428
rect 6015 60236 6032 60286
rect 6015 60094 6032 60144
rect 6015 59952 6032 60002
rect 6015 59810 6032 59860
rect 6015 59668 6032 59718
rect 6015 59526 6032 59576
rect 6015 59384 6032 59434
rect 6015 59242 6032 59292
rect 6015 59100 6032 59150
rect 6015 58958 6032 59008
rect 6015 58816 6032 58866
rect 6015 58674 6032 58724
rect 6015 58532 6032 58582
rect 6015 58390 6032 58440
rect 6015 58248 6032 58298
rect 6015 58106 6032 58156
rect 6015 57964 6032 58014
rect 6015 57822 6032 57872
rect 6015 57680 6032 57730
rect 6015 57538 6032 57588
rect 6015 57396 6032 57446
rect 6015 57254 6032 57304
rect 6015 57112 6032 57162
rect 6015 56970 6032 57020
rect 6015 56828 6032 56878
rect 6015 56686 6032 56736
rect 6015 56544 6032 56594
rect 6015 56402 6032 56452
rect 6015 56260 6032 56310
rect 6015 56118 6032 56168
rect 6015 55976 6032 56026
rect 6015 55834 6032 55884
rect 6015 55692 6032 55742
rect 6015 55550 6032 55600
rect 6015 55408 6032 55458
rect 6015 55266 6032 55316
rect 6015 55124 6032 55174
rect 6015 54982 6032 55032
rect 6015 54840 6032 54890
rect 6015 54698 6032 54748
rect 6015 54556 6032 54606
rect 6015 54414 6032 54464
rect 6015 54272 6032 54322
rect 6015 54130 6032 54180
rect 6015 53988 6032 54038
rect 6015 53846 6032 53896
rect 6015 53704 6032 53754
rect 6015 53562 6032 53612
rect 6015 53420 6032 53470
rect 6015 53278 6032 53328
rect 6015 53136 6032 53186
rect 6015 52994 6032 53044
rect 6015 52852 6032 52902
rect 6015 52710 6032 52760
rect 6015 52568 6032 52618
rect 6015 52426 6032 52476
rect 6015 52284 6032 52334
rect 6015 52142 6032 52192
rect 6015 52000 6032 52050
rect 6015 51858 6032 51908
rect 6015 51716 6032 51766
rect 6015 51574 6032 51624
rect 6015 51432 6032 51482
rect 6015 51290 6032 51340
rect 6015 51148 6032 51198
rect 6015 51006 6032 51056
rect 6015 50864 6032 50914
rect 6015 50722 6032 50772
rect 6015 50580 6032 50630
rect 6015 50438 6032 50488
rect 6015 50296 6032 50346
rect 6015 50154 6032 50204
rect 6015 50012 6032 50062
rect 6015 49870 6032 49920
rect 6015 49728 6032 49778
rect 6015 49586 6032 49636
rect 6015 49444 6032 49494
rect 6015 49302 6032 49352
rect 6015 49160 6032 49210
rect 6015 49018 6032 49068
rect 6015 48876 6032 48926
rect 6015 48734 6032 48784
rect 6015 48592 6032 48642
rect 6015 48450 6032 48500
rect 6015 48308 6032 48358
rect 6015 48166 6032 48216
rect 6015 48024 6032 48074
rect 6015 47882 6032 47932
rect 6015 47740 6032 47790
rect 6015 47598 6032 47648
rect 6015 47456 6032 47506
rect 6015 47314 6032 47364
rect 6015 47172 6032 47222
rect 6015 47030 6032 47080
rect 6015 46888 6032 46938
rect 6015 46746 6032 46796
rect 6015 46604 6032 46654
rect 6015 46462 6032 46512
rect 6015 46320 6032 46370
rect 6015 46178 6032 46228
rect 6015 46036 6032 46086
rect 6015 45894 6032 45944
rect 6015 45752 6032 45802
rect 6015 45610 6032 45660
rect 6015 45468 6032 45518
rect 6015 45326 6032 45376
rect 6015 45184 6032 45234
rect 6015 45042 6032 45092
rect 6015 44900 6032 44950
rect 6015 44758 6032 44808
rect 6015 44616 6032 44666
rect 6015 44474 6032 44524
rect 6015 44332 6032 44382
rect 6015 44190 6032 44240
rect 6015 44048 6032 44098
rect 6015 43906 6032 43956
rect 6015 43764 6032 43814
rect 6015 43622 6032 43672
rect 6015 43480 6032 43530
rect 6015 43338 6032 43388
rect 6015 43196 6032 43246
rect 6015 43054 6032 43104
rect 6015 42912 6032 42962
rect 6015 42770 6032 42820
rect 6015 42628 6032 42678
rect 6015 42486 6032 42536
rect 6015 42344 6032 42394
rect 6015 42202 6032 42252
rect 6015 42060 6032 42110
rect 6015 41918 6032 41968
rect 6015 41776 6032 41826
rect 6015 41634 6032 41684
rect 6015 41492 6032 41542
rect 6015 41350 6032 41400
rect 6015 41208 6032 41258
rect 6015 41066 6032 41116
rect 6015 40924 6032 40974
rect 6015 40782 6032 40832
rect 6015 40640 6032 40690
rect 6015 40498 6032 40548
rect 6015 40356 6032 40406
rect 6015 40214 6032 40264
rect 6015 40072 6032 40122
rect 6015 39930 6032 39980
rect 6015 39788 6032 39838
rect 6015 39646 6032 39696
rect 6015 39504 6032 39554
rect 6015 39362 6032 39412
rect 6015 39220 6032 39270
rect 6015 39078 6032 39128
rect 6015 38936 6032 38986
rect 6015 38794 6032 38844
rect 6015 38652 6032 38702
rect 6015 38510 6032 38560
rect 6015 38368 6032 38418
rect 6015 38226 6032 38276
rect 6015 38084 6032 38134
rect 6015 37942 6032 37992
rect 6015 37800 6032 37850
rect 6015 37658 6032 37708
rect 6015 37516 6032 37566
rect 6015 37374 6032 37424
rect 6015 37232 6032 37282
rect 6015 37090 6032 37140
rect 6015 36948 6032 36998
rect 6015 36806 6032 36856
rect 6015 36664 6032 36714
rect 6015 36522 6032 36572
rect 6015 36380 6032 36430
rect 6015 36238 6032 36288
rect 6015 36096 6032 36146
rect 6015 35954 6032 36004
rect 6015 35812 6032 35862
rect 6015 35670 6032 35720
rect 6015 35528 6032 35578
rect 6015 35386 6032 35436
rect 6015 35244 6032 35294
rect 6015 35102 6032 35152
rect 6015 34960 6032 35010
rect 6015 34818 6032 34868
rect 6015 34676 6032 34726
rect 6015 34534 6032 34584
rect 6015 34392 6032 34442
rect 6015 34250 6032 34300
rect 6015 34108 6032 34158
rect 6015 33966 6032 34016
rect 6015 33824 6032 33874
rect 6015 33682 6032 33732
rect 6015 33540 6032 33590
rect 6015 33398 6032 33448
rect 6015 33256 6032 33306
rect 6015 33114 6032 33164
rect 6015 32972 6032 33022
rect 6015 32830 6032 32880
rect 6015 32688 6032 32738
rect 6015 32546 6032 32596
rect 6015 32404 6032 32454
rect 6015 32262 6032 32312
rect 6015 32120 6032 32170
rect 6015 31978 6032 32028
rect 6015 31836 6032 31886
rect 6015 31694 6032 31744
rect 6015 31552 6032 31602
rect 6015 31410 6032 31460
rect 6015 31268 6032 31318
rect 6015 31126 6032 31176
rect 6015 30984 6032 31034
rect 6015 30842 6032 30892
rect 6015 30700 6032 30750
rect 6015 30558 6032 30608
rect 6015 30416 6032 30466
rect 6015 30274 6032 30324
rect 6015 30132 6032 30182
rect 6015 29990 6032 30040
rect 6015 29848 6032 29898
rect 6015 29706 6032 29756
rect 6015 29564 6032 29614
rect 6015 29422 6032 29472
rect 6015 29280 6032 29330
rect 6015 29138 6032 29188
rect 6015 28996 6032 29046
rect 6015 28854 6032 28904
rect 6015 28712 6032 28762
rect 6015 28570 6032 28620
rect 6015 28428 6032 28478
rect 6015 28286 6032 28336
rect 6015 28144 6032 28194
rect 6015 28002 6032 28052
rect 6015 27860 6032 27910
rect 6015 27718 6032 27768
rect 6015 27576 6032 27626
rect 6015 27434 6032 27484
rect 6015 27292 6032 27342
rect 6015 27150 6032 27200
rect 6015 27008 6032 27058
rect 6015 26866 6032 26916
rect 6015 26724 6032 26774
rect 6015 26582 6032 26632
rect 6015 26440 6032 26490
rect 6015 26298 6032 26348
rect 6015 26156 6032 26206
rect 6015 26014 6032 26064
rect 6015 25872 6032 25922
rect 6015 25730 6032 25780
rect 6015 25588 6032 25638
rect 6015 25446 6032 25496
rect 6015 25304 6032 25354
rect 6015 25162 6032 25212
rect 6015 25020 6032 25070
rect 6015 24878 6032 24928
rect 6015 24736 6032 24786
rect 6015 24594 6032 24644
rect 6015 24452 6032 24502
rect 6015 24310 6032 24360
rect 6015 24168 6032 24218
rect 6015 24026 6032 24076
rect 6015 23884 6032 23934
rect 6015 23742 6032 23792
rect 6015 23600 6032 23650
rect 6015 23458 6032 23508
rect 6015 23316 6032 23366
rect 6015 23174 6032 23224
rect 6015 23032 6032 23082
rect 6015 22890 6032 22940
rect 6015 22748 6032 22798
rect 6015 22606 6032 22656
rect 6015 22464 6032 22514
rect 6015 22322 6032 22372
rect 6015 22180 6032 22230
rect 6015 22038 6032 22088
rect 6015 21896 6032 21946
rect 6015 21754 6032 21804
rect 6015 21612 6032 21662
rect 6015 21470 6032 21520
rect 6015 21328 6032 21378
rect 6015 21186 6032 21236
rect 6015 21044 6032 21094
rect 6015 20902 6032 20952
rect 6015 20760 6032 20810
rect 6015 20618 6032 20668
rect 6015 20476 6032 20526
rect 6015 20334 6032 20384
rect 6015 20192 6032 20242
rect 6015 20050 6032 20100
rect 6015 19908 6032 19958
rect 6015 19766 6032 19816
rect 6015 19624 6032 19674
rect 6015 19482 6032 19532
rect 6015 19340 6032 19390
rect 6015 19198 6032 19248
rect 6015 19056 6032 19106
rect 6015 18914 6032 18964
rect 6015 18772 6032 18822
rect 6015 18630 6032 18680
rect 6015 18488 6032 18538
rect 6015 18346 6032 18396
rect 6015 18204 6032 18254
rect 6015 18062 6032 18112
rect 6015 17920 6032 17970
rect 6015 17778 6032 17828
rect 6015 17636 6032 17686
rect 6015 17494 6032 17544
rect 6015 17352 6032 17402
rect 6015 17210 6032 17260
rect 6015 17068 6032 17118
rect 6015 16926 6032 16976
rect 6015 16784 6032 16834
rect 6015 16642 6032 16692
rect 6015 16500 6032 16550
rect 6015 16358 6032 16408
rect 6015 16216 6032 16266
rect 6015 16074 6032 16124
rect 6015 15932 6032 15982
rect 6015 15790 6032 15840
rect 6015 15648 6032 15698
rect 6015 15506 6032 15556
rect 6015 15364 6032 15414
rect 6015 15222 6032 15272
rect 6015 15080 6032 15130
rect 6015 14938 6032 14988
rect 6015 14796 6032 14846
rect 6015 14654 6032 14704
rect 6015 14512 6032 14562
rect 6015 14370 6032 14420
rect 6015 14228 6032 14278
rect 6015 14086 6032 14136
rect 6015 13944 6032 13994
rect 6015 13802 6032 13852
rect 6015 13660 6032 13710
rect 6015 13518 6032 13568
rect 6015 13376 6032 13426
rect 6015 13234 6032 13284
rect 6015 13092 6032 13142
rect 6015 12950 6032 13000
rect 6015 12808 6032 12858
rect 6015 12666 6032 12716
rect 6015 12524 6032 12574
rect 6015 12382 6032 12432
rect 6015 12240 6032 12290
rect 6015 12098 6032 12148
rect 6015 11956 6032 12006
rect 6015 11814 6032 11864
rect 6015 11672 6032 11722
rect 6015 11530 6032 11580
rect 6015 11388 6032 11438
rect 6015 11246 6032 11296
rect 6015 11104 6032 11154
rect 6015 10962 6032 11012
rect 6015 10820 6032 10870
rect 6015 10678 6032 10728
rect 6015 10536 6032 10586
rect 6015 10394 6032 10444
rect 6015 10252 6032 10302
rect 6015 10110 6032 10160
rect 6015 9968 6032 10018
rect 6015 9826 6032 9876
rect 6015 9684 6032 9734
rect 6015 9542 6032 9592
rect 6015 9400 6032 9450
rect 6015 9258 6032 9308
rect 6015 9116 6032 9166
rect 6015 8974 6032 9024
rect 6015 8832 6032 8882
rect 6015 8690 6032 8740
rect 6015 8548 6032 8598
rect 6015 8406 6032 8456
rect 6015 8264 6032 8314
rect 6015 8122 6032 8172
rect 6015 7980 6032 8030
rect 6015 7838 6032 7888
rect 6015 7696 6032 7746
rect 6015 7554 6032 7604
rect 6015 7412 6032 7462
rect 6015 7270 6032 7320
rect 6015 7128 6032 7178
rect 6015 6986 6032 7036
rect 6015 6844 6032 6894
rect 6015 6702 6032 6752
rect 6015 6560 6032 6610
rect 6015 6418 6032 6468
rect 6015 6276 6032 6326
rect 6015 6134 6032 6184
rect 6015 5992 6032 6042
rect 6015 5850 6032 5900
rect 6015 5708 6032 5758
rect 6015 5566 6032 5616
rect 6015 5424 6032 5474
rect 6015 5282 6032 5332
rect 6015 5140 6032 5190
rect 6015 4998 6032 5048
rect 6015 4856 6032 4906
rect 6015 4714 6032 4764
rect 6015 4572 6032 4622
rect 6015 4430 6032 4480
rect 6015 4288 6032 4338
rect 6015 4146 6032 4196
rect 6015 4004 6032 4054
rect 6015 3862 6032 3912
rect 6015 3720 6032 3770
rect 6015 3578 6032 3628
rect 6015 3436 6032 3486
rect 6015 3294 6032 3344
rect 6015 3152 6032 3202
rect 6015 3010 6032 3060
rect 6015 2868 6032 2918
rect 6015 2726 6032 2776
rect 6015 2584 6032 2634
rect 6015 2442 6032 2492
rect 6015 2300 6032 2350
rect 6015 2158 6032 2208
rect 6015 2016 6032 2066
rect 6015 1874 6032 1924
rect 6015 1732 6032 1782
rect 6015 1590 6032 1640
rect 6015 1448 6032 1498
rect 6015 1306 6032 1356
rect 6015 1164 6032 1214
rect 6015 1022 6032 1072
rect 6015 880 6032 930
rect 6015 738 6032 788
rect 6015 596 6032 646
rect 6015 454 6032 504
rect 6015 312 6032 362
rect 6015 170 6032 220
rect 56 -128 100 -84
rect 6108 6 6174 60
rect 6440 9 6506 75
rect 6606 7 6672 73
rect 6938 13 7004 67
rect 7104 6 7170 60
rect 7436 6 7502 72
rect 7602 6 7668 60
rect 7934 9 8000 75
rect 5554 -134 5598 -78
rect 5733 -713 5787 -659
rect 6039 -715 6093 -661
rect 6341 -715 6395 -661
rect 6653 -713 6707 -659
rect 6967 -717 7021 -663
rect 7263 -723 7317 -669
rect 7565 -715 7619 -661
rect 7883 -715 7937 -661
<< metal1 >>
rect 5978 146048 6034 146060
rect 5752 146042 5984 146048
rect 5752 145998 5764 146042
rect 5808 145998 5984 146042
rect 5752 145992 5984 145998
rect 6028 145992 6034 146048
rect 5978 145980 6034 145992
rect -974 145860 -926 145866
rect -974 145854 96 145860
rect -974 145818 -968 145854
rect -932 145818 36 145854
rect 84 145818 96 145854
rect -974 145812 96 145818
rect -974 145806 -926 145812
rect 5714 145486 6040 145504
rect 5714 145436 6015 145486
rect 6032 145436 6040 145486
rect 5714 145418 6040 145436
rect 5714 145344 6040 145362
rect 5714 145294 6015 145344
rect 6032 145294 6040 145344
rect -232 145276 -152 145286
rect 5714 145276 6040 145294
rect -232 145220 -222 145276
rect -164 145220 -152 145276
rect -232 145210 -152 145220
rect 5714 145202 6040 145220
rect 5714 145152 6015 145202
rect 6032 145152 6040 145202
rect 5714 145134 6040 145152
rect 5714 145060 6040 145078
rect 5714 145010 6015 145060
rect 6032 145010 6040 145060
rect 5714 144992 6040 145010
rect 5714 144918 6040 144936
rect 5714 144868 6015 144918
rect 6032 144868 6040 144918
rect 5714 144850 6040 144868
rect 5714 144776 6040 144794
rect 5714 144726 6015 144776
rect 6032 144726 6040 144776
rect 5714 144708 6040 144726
rect 5714 144634 6040 144652
rect 5714 144584 6015 144634
rect 6032 144584 6040 144634
rect 5714 144566 6040 144584
rect 5714 144492 6040 144510
rect 5714 144442 6015 144492
rect 6032 144442 6040 144492
rect 5714 144424 6040 144442
rect 5714 144350 6040 144368
rect 5714 144300 6015 144350
rect 6032 144300 6040 144350
rect 5714 144282 6040 144300
rect 5714 144208 6040 144226
rect 5714 144158 6015 144208
rect 6032 144158 6040 144208
rect 5714 144140 6040 144158
rect 5714 144066 6040 144084
rect 5714 144016 6015 144066
rect 6032 144016 6040 144066
rect 5714 143998 6040 144016
rect 5714 143924 6040 143942
rect 5714 143874 6015 143924
rect 6032 143874 6040 143924
rect 5714 143856 6040 143874
rect 5714 143782 6040 143800
rect 5714 143732 6015 143782
rect 6032 143732 6040 143782
rect 5714 143714 6040 143732
rect 5714 143640 6040 143658
rect 5714 143590 6015 143640
rect 6032 143590 6040 143640
rect 5714 143572 6040 143590
rect 5714 143498 6040 143516
rect 5714 143448 6015 143498
rect 6032 143448 6040 143498
rect 5714 143430 6040 143448
rect 5714 143356 6040 143374
rect 5714 143306 6015 143356
rect 6032 143306 6040 143356
rect 5714 143288 6040 143306
rect 5714 143214 6040 143232
rect 5714 143164 6015 143214
rect 6032 143164 6040 143214
rect 5714 143146 6040 143164
rect 5714 143072 6040 143090
rect 5714 143022 6015 143072
rect 6032 143022 6040 143072
rect 5714 143004 6040 143022
rect 5714 142930 6040 142948
rect 5714 142880 6015 142930
rect 6032 142880 6040 142930
rect 5714 142862 6040 142880
rect 5714 142788 6040 142806
rect 5714 142738 6015 142788
rect 6032 142738 6040 142788
rect 5714 142720 6040 142738
rect 5714 142646 6040 142664
rect 5714 142596 6015 142646
rect 6032 142596 6040 142646
rect 5714 142578 6040 142596
rect 5714 142504 6040 142522
rect 5714 142454 6015 142504
rect 6032 142454 6040 142504
rect 5714 142436 6040 142454
rect -172 142385 -86 142396
rect -401 142319 -161 142385
rect -95 142319 -86 142385
rect -172 142310 -86 142319
rect 5714 142362 6040 142380
rect 5714 142312 6015 142362
rect 6032 142312 6040 142362
rect 5714 142294 6040 142312
rect 5714 142220 6040 142238
rect 5714 142170 6015 142220
rect 6032 142170 6040 142220
rect 5714 142152 6040 142170
rect 5714 142078 6040 142096
rect 5714 142028 6015 142078
rect 6032 142028 6040 142078
rect 5714 142010 6040 142028
rect 5714 141936 6040 141954
rect 5714 141886 6015 141936
rect 6032 141886 6040 141936
rect 5714 141868 6040 141886
rect 5714 141794 6040 141812
rect 5714 141744 6015 141794
rect 6032 141744 6040 141794
rect 5714 141726 6040 141744
rect 5714 141652 6040 141670
rect 5714 141602 6015 141652
rect 6032 141602 6040 141652
rect 5714 141584 6040 141602
rect 5714 141510 6040 141528
rect 5714 141460 6015 141510
rect 6032 141460 6040 141510
rect 5714 141442 6040 141460
rect 5714 141368 6040 141386
rect 5714 141318 6015 141368
rect 6032 141318 6040 141368
rect 5714 141300 6040 141318
rect 5714 141226 6040 141244
rect 5714 141176 6015 141226
rect 6032 141176 6040 141226
rect 5714 141158 6040 141176
rect 5714 141084 6040 141102
rect 5714 141034 6015 141084
rect 6032 141034 6040 141084
rect 5714 141016 6040 141034
rect 5714 140942 6040 140960
rect 5714 140892 6015 140942
rect 6032 140892 6040 140942
rect 5714 140874 6040 140892
rect 5714 140800 6040 140818
rect 5714 140750 6015 140800
rect 6032 140750 6040 140800
rect 5714 140732 6040 140750
rect 5714 140658 6040 140676
rect 5714 140608 6015 140658
rect 6032 140608 6040 140658
rect 5714 140590 6040 140608
rect 5714 140516 6040 140534
rect 5714 140466 6015 140516
rect 6032 140466 6040 140516
rect 5714 140448 6040 140466
rect 5714 140374 6040 140392
rect 5714 140324 6015 140374
rect 6032 140324 6040 140374
rect 5714 140306 6040 140324
rect 5714 140232 6040 140250
rect 5714 140182 6015 140232
rect 6032 140182 6040 140232
rect 5714 140164 6040 140182
rect 5714 140090 6040 140108
rect 5714 140040 6015 140090
rect 6032 140040 6040 140090
rect 5714 140022 6040 140040
rect 5714 139948 6040 139966
rect 5714 139898 6015 139948
rect 6032 139898 6040 139948
rect 5714 139880 6040 139898
rect 5714 139806 6040 139824
rect 5714 139756 6015 139806
rect 6032 139756 6040 139806
rect 5714 139738 6040 139756
rect 5714 139664 6040 139682
rect 5714 139614 6015 139664
rect 6032 139614 6040 139664
rect 5714 139596 6040 139614
rect 5714 139522 6040 139540
rect 5714 139472 6015 139522
rect 6032 139472 6040 139522
rect 5714 139454 6040 139472
rect 5714 139380 6040 139398
rect 5714 139330 6015 139380
rect 6032 139330 6040 139380
rect 5714 139312 6040 139330
rect 5714 139238 6040 139256
rect 5714 139188 6015 139238
rect 6032 139188 6040 139238
rect 5714 139170 6040 139188
rect -182 139130 -104 139138
rect -399 139064 -177 139130
rect -111 139064 -104 139130
rect -182 139058 -104 139064
rect 5714 139096 6040 139114
rect 5714 139046 6015 139096
rect 6032 139046 6040 139096
rect 5714 139028 6040 139046
rect 5714 138954 6040 138972
rect 5714 138904 6015 138954
rect 6032 138904 6040 138954
rect 5714 138886 6040 138904
rect 5714 138812 6040 138830
rect 5714 138762 6015 138812
rect 6032 138762 6040 138812
rect 5714 138744 6040 138762
rect 5714 138670 6040 138688
rect 5714 138620 6015 138670
rect 6032 138620 6040 138670
rect 5714 138602 6040 138620
rect 5714 138528 6040 138546
rect 5714 138478 6015 138528
rect 6032 138478 6040 138528
rect 5714 138460 6040 138478
rect 5714 138386 6040 138404
rect 5714 138336 6015 138386
rect 6032 138336 6040 138386
rect 5714 138318 6040 138336
rect 5714 138244 6040 138262
rect 5714 138194 6015 138244
rect 6032 138194 6040 138244
rect 5714 138176 6040 138194
rect 5714 138102 6040 138120
rect 5714 138052 6015 138102
rect 6032 138052 6040 138102
rect 5714 138034 6040 138052
rect 5714 137960 6040 137978
rect 5714 137910 6015 137960
rect 6032 137910 6040 137960
rect 5714 137892 6040 137910
rect 5714 137818 6040 137836
rect 5714 137768 6015 137818
rect 6032 137768 6040 137818
rect 5714 137750 6040 137768
rect 5714 137676 6040 137694
rect 5714 137626 6015 137676
rect 6032 137626 6040 137676
rect 5714 137608 6040 137626
rect 5714 137534 6040 137552
rect 5714 137484 6015 137534
rect 6032 137484 6040 137534
rect 5714 137466 6040 137484
rect 5714 137392 6040 137410
rect 5714 137342 6015 137392
rect 6032 137342 6040 137392
rect 5714 137324 6040 137342
rect 5714 137250 6040 137268
rect 5714 137200 6015 137250
rect 6032 137200 6040 137250
rect 5714 137182 6040 137200
rect 5714 137108 6040 137126
rect 5714 137058 6015 137108
rect 6032 137058 6040 137108
rect 5714 137040 6040 137058
rect 5714 136966 6040 136984
rect 5714 136916 6015 136966
rect 6032 136916 6040 136966
rect 5714 136898 6040 136916
rect 5714 136824 6040 136842
rect 5714 136774 6015 136824
rect 6032 136774 6040 136824
rect 5714 136756 6040 136774
rect 5714 136682 6040 136700
rect 5714 136632 6015 136682
rect 6032 136632 6040 136682
rect 5714 136614 6040 136632
rect 5714 136540 6040 136558
rect 5714 136490 6015 136540
rect 6032 136490 6040 136540
rect 5714 136472 6040 136490
rect 5714 136398 6040 136416
rect 5714 136348 6015 136398
rect 6032 136348 6040 136398
rect 5714 136330 6040 136348
rect 5714 136256 6040 136274
rect 5714 136206 6015 136256
rect 6032 136206 6040 136256
rect 5714 136188 6040 136206
rect 5714 136114 6040 136132
rect 5714 136064 6015 136114
rect 6032 136064 6040 136114
rect 5714 136046 6040 136064
rect 5714 135972 6040 135990
rect -150 135919 -74 135932
rect -150 135917 -138 135919
rect -392 135868 -138 135917
rect -150 135867 -138 135868
rect -86 135867 -74 135919
rect 5714 135922 6015 135972
rect 6032 135922 6040 135972
rect 5714 135904 6040 135922
rect -150 135856 -74 135867
rect 5714 135830 6040 135848
rect 5714 135780 6015 135830
rect 6032 135780 6040 135830
rect 5714 135762 6040 135780
rect 5714 135688 6040 135706
rect 5714 135638 6015 135688
rect 6032 135638 6040 135688
rect 5714 135620 6040 135638
rect 5714 135546 6040 135564
rect 5714 135496 6015 135546
rect 6032 135496 6040 135546
rect 5714 135478 6040 135496
rect 5714 135404 6040 135422
rect 5714 135354 6015 135404
rect 6032 135354 6040 135404
rect 5714 135336 6040 135354
rect 5714 135262 6040 135280
rect 5714 135212 6015 135262
rect 6032 135212 6040 135262
rect 5714 135194 6040 135212
rect 5714 135120 6040 135138
rect 5714 135070 6015 135120
rect 6032 135070 6040 135120
rect 5714 135052 6040 135070
rect 5714 134978 6040 134996
rect 5714 134928 6015 134978
rect 6032 134928 6040 134978
rect 5714 134910 6040 134928
rect 5714 134836 6040 134854
rect 5714 134786 6015 134836
rect 6032 134786 6040 134836
rect 5714 134768 6040 134786
rect 5714 134694 6040 134712
rect 5714 134644 6015 134694
rect 6032 134644 6040 134694
rect 5714 134626 6040 134644
rect 5714 134552 6040 134570
rect 5714 134502 6015 134552
rect 6032 134502 6040 134552
rect 5714 134484 6040 134502
rect 5714 134410 6040 134428
rect 5714 134360 6015 134410
rect 6032 134360 6040 134410
rect 5714 134342 6040 134360
rect 5714 134268 6040 134286
rect 5714 134218 6015 134268
rect 6032 134218 6040 134268
rect 5714 134200 6040 134218
rect 5714 134126 6040 134144
rect 5714 134076 6015 134126
rect 6032 134076 6040 134126
rect 5714 134058 6040 134076
rect 5714 133984 6040 134002
rect 5714 133934 6015 133984
rect 6032 133934 6040 133984
rect 5714 133916 6040 133934
rect 5714 133842 6040 133860
rect 5714 133792 6015 133842
rect 6032 133792 6040 133842
rect 5714 133774 6040 133792
rect 5714 133700 6040 133718
rect 5714 133650 6015 133700
rect 6032 133650 6040 133700
rect 5714 133632 6040 133650
rect 5714 133558 6040 133576
rect 5714 133508 6015 133558
rect 6032 133508 6040 133558
rect 5714 133490 6040 133508
rect 5714 133416 6040 133434
rect 5714 133366 6015 133416
rect 6032 133366 6040 133416
rect 5714 133348 6040 133366
rect 5714 133274 6040 133292
rect 5714 133224 6015 133274
rect 6032 133224 6040 133274
rect 5714 133206 6040 133224
rect 5714 133132 6040 133150
rect 5714 133082 6015 133132
rect 6032 133082 6040 133132
rect 5714 133064 6040 133082
rect 5714 132990 6040 133008
rect 5714 132940 6015 132990
rect 6032 132940 6040 132990
rect 5714 132922 6040 132940
rect 5714 132848 6040 132866
rect 5714 132798 6015 132848
rect 6032 132798 6040 132848
rect 5714 132780 6040 132798
rect 5714 132706 6040 132724
rect -144 132659 -60 132668
rect -401 132593 -135 132659
rect -69 132593 -60 132659
rect 5714 132656 6015 132706
rect 6032 132656 6040 132706
rect 5714 132638 6040 132656
rect -144 132582 -60 132593
rect 5714 132564 6040 132582
rect 5714 132514 6015 132564
rect 6032 132514 6040 132564
rect 5714 132496 6040 132514
rect 5714 132422 6040 132440
rect 5714 132372 6015 132422
rect 6032 132372 6040 132422
rect 5714 132354 6040 132372
rect 5714 132280 6040 132298
rect 5714 132230 6015 132280
rect 6032 132230 6040 132280
rect 5714 132212 6040 132230
rect 5714 132138 6040 132156
rect 5714 132088 6015 132138
rect 6032 132088 6040 132138
rect 5714 132070 6040 132088
rect 5714 131996 6040 132014
rect 5714 131946 6015 131996
rect 6032 131946 6040 131996
rect 5714 131928 6040 131946
rect 5714 131854 6040 131872
rect 5714 131804 6015 131854
rect 6032 131804 6040 131854
rect 5714 131786 6040 131804
rect 5714 131712 6040 131730
rect 5714 131662 6015 131712
rect 6032 131662 6040 131712
rect 5714 131644 6040 131662
rect 5714 131570 6040 131588
rect 5714 131520 6015 131570
rect 6032 131520 6040 131570
rect 5714 131502 6040 131520
rect 5714 131428 6040 131446
rect 5714 131378 6015 131428
rect 6032 131378 6040 131428
rect 5714 131360 6040 131378
rect 5714 131286 6040 131304
rect 5714 131236 6015 131286
rect 6032 131236 6040 131286
rect 5714 131218 6040 131236
rect 5714 131144 6040 131162
rect 5714 131094 6015 131144
rect 6032 131094 6040 131144
rect 5714 131076 6040 131094
rect 5714 131002 6040 131020
rect 5714 130952 6015 131002
rect 6032 130952 6040 131002
rect 5714 130934 6040 130952
rect 5714 130860 6040 130878
rect 5714 130810 6015 130860
rect 6032 130810 6040 130860
rect 5714 130792 6040 130810
rect 5714 130718 6040 130736
rect 5714 130668 6015 130718
rect 6032 130668 6040 130718
rect 5714 130650 6040 130668
rect 5714 130576 6040 130594
rect 5714 130526 6015 130576
rect 6032 130526 6040 130576
rect 5714 130508 6040 130526
rect 5714 130434 6040 130452
rect 5714 130384 6015 130434
rect 6032 130384 6040 130434
rect 5714 130366 6040 130384
rect 5714 130292 6040 130310
rect 5714 130242 6015 130292
rect 6032 130242 6040 130292
rect 5714 130224 6040 130242
rect 5714 130150 6040 130168
rect 5714 130100 6015 130150
rect 6032 130100 6040 130150
rect 5714 130082 6040 130100
rect 5714 130008 6040 130026
rect 5714 129958 6015 130008
rect 6032 129958 6040 130008
rect 5714 129940 6040 129958
rect 5714 129866 6040 129884
rect 5714 129816 6015 129866
rect 6032 129816 6040 129866
rect 5714 129798 6040 129816
rect 5714 129724 6040 129742
rect 5714 129674 6015 129724
rect 6032 129674 6040 129724
rect 5714 129656 6040 129674
rect 5714 129582 6040 129600
rect 5714 129532 6015 129582
rect 6032 129532 6040 129582
rect 5714 129514 6040 129532
rect 5714 129440 6040 129458
rect -128 129425 -44 129434
rect -401 129359 -119 129425
rect -53 129359 -44 129425
rect 5714 129390 6015 129440
rect 6032 129390 6040 129440
rect 5714 129372 6040 129390
rect -128 129350 -44 129359
rect 5714 129298 6040 129316
rect 5714 129248 6015 129298
rect 6032 129248 6040 129298
rect 5714 129230 6040 129248
rect 5714 129156 6040 129174
rect 5714 129106 6015 129156
rect 6032 129106 6040 129156
rect 5714 129088 6040 129106
rect 5714 129014 6040 129032
rect 5714 128964 6015 129014
rect 6032 128964 6040 129014
rect 5714 128946 6040 128964
rect 5714 128872 6040 128890
rect 5714 128822 6015 128872
rect 6032 128822 6040 128872
rect 5714 128804 6040 128822
rect 5714 128730 6040 128748
rect 5714 128680 6015 128730
rect 6032 128680 6040 128730
rect 5714 128662 6040 128680
rect 5714 128588 6040 128606
rect 5714 128538 6015 128588
rect 6032 128538 6040 128588
rect 5714 128520 6040 128538
rect 5714 128446 6040 128464
rect 5714 128396 6015 128446
rect 6032 128396 6040 128446
rect 5714 128378 6040 128396
rect 5714 128304 6040 128322
rect 5714 128254 6015 128304
rect 6032 128254 6040 128304
rect 5714 128236 6040 128254
rect 5714 128162 6040 128180
rect 5714 128112 6015 128162
rect 6032 128112 6040 128162
rect 5714 128094 6040 128112
rect 5714 128020 6040 128038
rect 5714 127970 6015 128020
rect 6032 127970 6040 128020
rect 5714 127952 6040 127970
rect 5714 127878 6040 127896
rect 5714 127828 6015 127878
rect 6032 127828 6040 127878
rect 5714 127810 6040 127828
rect 5714 127736 6040 127754
rect 5714 127686 6015 127736
rect 6032 127686 6040 127736
rect 5714 127668 6040 127686
rect 5714 127594 6040 127612
rect 5714 127544 6015 127594
rect 6032 127544 6040 127594
rect 5714 127526 6040 127544
rect 5714 127452 6040 127470
rect 5714 127402 6015 127452
rect 6032 127402 6040 127452
rect 5714 127384 6040 127402
rect 5714 127310 6040 127328
rect 5714 127260 6015 127310
rect 6032 127260 6040 127310
rect 5714 127242 6040 127260
rect 5714 127168 6040 127186
rect 5714 127118 6015 127168
rect 6032 127118 6040 127168
rect 5714 127100 6040 127118
rect 5714 127026 6040 127044
rect 5714 126976 6015 127026
rect 6032 126976 6040 127026
rect 5714 126958 6040 126976
rect 5714 126884 6040 126902
rect 5714 126834 6015 126884
rect 6032 126834 6040 126884
rect 5714 126816 6040 126834
rect 5714 126742 6040 126760
rect 5714 126692 6015 126742
rect 6032 126692 6040 126742
rect 5714 126674 6040 126692
rect 5714 126600 6040 126618
rect 5714 126550 6015 126600
rect 6032 126550 6040 126600
rect 5714 126532 6040 126550
rect 5714 126458 6040 126476
rect 5714 126408 6015 126458
rect 6032 126408 6040 126458
rect 5714 126390 6040 126408
rect 5714 126316 6040 126334
rect 5714 126266 6015 126316
rect 6032 126266 6040 126316
rect 5714 126248 6040 126266
rect -144 126183 -60 126192
rect -401 126117 -139 126183
rect -73 126117 -60 126183
rect -144 126108 -60 126117
rect 5714 126174 6040 126192
rect 5714 126124 6015 126174
rect 6032 126124 6040 126174
rect 5714 126106 6040 126124
rect 5714 126032 6040 126050
rect 5714 125982 6015 126032
rect 6032 125982 6040 126032
rect 5714 125964 6040 125982
rect 5714 125890 6040 125908
rect 5714 125840 6015 125890
rect 6032 125840 6040 125890
rect 5714 125822 6040 125840
rect 5714 125748 6040 125766
rect 5714 125698 6015 125748
rect 6032 125698 6040 125748
rect 5714 125680 6040 125698
rect 5714 125606 6040 125624
rect 5714 125556 6015 125606
rect 6032 125556 6040 125606
rect 5714 125538 6040 125556
rect 5714 125464 6040 125482
rect 5714 125414 6015 125464
rect 6032 125414 6040 125464
rect 5714 125396 6040 125414
rect 5714 125322 6040 125340
rect 5714 125272 6015 125322
rect 6032 125272 6040 125322
rect 5714 125254 6040 125272
rect 5714 125180 6040 125198
rect 5714 125130 6015 125180
rect 6032 125130 6040 125180
rect 5714 125112 6040 125130
rect 5714 125038 6040 125056
rect 5714 124988 6015 125038
rect 6032 124988 6040 125038
rect 5714 124970 6040 124988
rect 5714 124896 6040 124914
rect 5714 124846 6015 124896
rect 6032 124846 6040 124896
rect 5714 124828 6040 124846
rect 5714 124754 6040 124772
rect 5714 124704 6015 124754
rect 6032 124704 6040 124754
rect 5714 124686 6040 124704
rect 5714 124612 6040 124630
rect 5714 124562 6015 124612
rect 6032 124562 6040 124612
rect 5714 124544 6040 124562
rect 5714 124470 6040 124488
rect 5714 124420 6015 124470
rect 6032 124420 6040 124470
rect 5714 124402 6040 124420
rect 5714 124328 6040 124346
rect 5714 124278 6015 124328
rect 6032 124278 6040 124328
rect 5714 124260 6040 124278
rect 5714 124186 6040 124204
rect 5714 124136 6015 124186
rect 6032 124136 6040 124186
rect 5714 124118 6040 124136
rect 5714 124044 6040 124062
rect 5714 123994 6015 124044
rect 6032 123994 6040 124044
rect 5714 123976 6040 123994
rect 5714 123902 6040 123920
rect 5714 123852 6015 123902
rect 6032 123852 6040 123902
rect 5714 123834 6040 123852
rect 5714 123760 6040 123778
rect 5714 123710 6015 123760
rect 6032 123710 6040 123760
rect 5714 123692 6040 123710
rect 5714 123618 6040 123636
rect 5714 123568 6015 123618
rect 6032 123568 6040 123618
rect 5714 123550 6040 123568
rect 5714 123476 6040 123494
rect 5714 123426 6015 123476
rect 6032 123426 6040 123476
rect 5714 123408 6040 123426
rect 5714 123334 6040 123352
rect 5714 123284 6015 123334
rect 6032 123284 6040 123334
rect 5714 123266 6040 123284
rect 5714 123192 6040 123210
rect 5714 123142 6015 123192
rect 6032 123142 6040 123192
rect 5714 123124 6040 123142
rect 5714 123050 6040 123068
rect 5714 123000 6015 123050
rect 6032 123000 6040 123050
rect 5714 122982 6040 123000
rect -166 122951 -82 122960
rect -401 122885 -157 122951
rect -91 122885 -82 122951
rect -166 122876 -82 122885
rect 5714 122908 6040 122926
rect 5714 122858 6015 122908
rect 6032 122858 6040 122908
rect 5714 122840 6040 122858
rect 5714 122766 6040 122784
rect 5714 122716 6015 122766
rect 6032 122716 6040 122766
rect 5714 122698 6040 122716
rect 5714 122624 6040 122642
rect 5714 122574 6015 122624
rect 6032 122574 6040 122624
rect 5714 122556 6040 122574
rect 5714 122482 6040 122500
rect 5714 122432 6015 122482
rect 6032 122432 6040 122482
rect 5714 122414 6040 122432
rect 5714 122340 6040 122358
rect 5714 122290 6015 122340
rect 6032 122290 6040 122340
rect 5714 122272 6040 122290
rect 5714 122198 6040 122216
rect 5714 122148 6015 122198
rect 6032 122148 6040 122198
rect 5714 122130 6040 122148
rect 5714 122056 6040 122074
rect 5714 122006 6015 122056
rect 6032 122006 6040 122056
rect 5714 121988 6040 122006
rect 5714 121914 6040 121932
rect 5714 121864 6015 121914
rect 6032 121864 6040 121914
rect 5714 121846 6040 121864
rect 5714 121772 6040 121790
rect 5714 121722 6015 121772
rect 6032 121722 6040 121772
rect 5714 121704 6040 121722
rect 5714 121630 6040 121648
rect 5714 121580 6015 121630
rect 6032 121580 6040 121630
rect 5714 121562 6040 121580
rect 5714 121488 6040 121506
rect 5714 121438 6015 121488
rect 6032 121438 6040 121488
rect 5714 121420 6040 121438
rect 5714 121346 6040 121364
rect 5714 121296 6015 121346
rect 6032 121296 6040 121346
rect 5714 121278 6040 121296
rect 5714 121204 6040 121222
rect 5714 121154 6015 121204
rect 6032 121154 6040 121204
rect 5714 121136 6040 121154
rect 5714 121062 6040 121080
rect 5714 121012 6015 121062
rect 6032 121012 6040 121062
rect 5714 120994 6040 121012
rect 5714 120920 6040 120938
rect 5714 120870 6015 120920
rect 6032 120870 6040 120920
rect 5714 120852 6040 120870
rect 5714 120778 6040 120796
rect 5714 120728 6015 120778
rect 6032 120728 6040 120778
rect 5714 120710 6040 120728
rect 5714 120636 6040 120654
rect 5714 120586 6015 120636
rect 6032 120586 6040 120636
rect 5714 120568 6040 120586
rect 5714 120494 6040 120512
rect 5714 120444 6015 120494
rect 6032 120444 6040 120494
rect 5714 120426 6040 120444
rect 5714 120352 6040 120370
rect 5714 120302 6015 120352
rect 6032 120302 6040 120352
rect 5714 120284 6040 120302
rect 5714 120210 6040 120228
rect 5714 120160 6015 120210
rect 6032 120160 6040 120210
rect 5714 120142 6040 120160
rect 5714 120068 6040 120086
rect 5714 120018 6015 120068
rect 6032 120018 6040 120068
rect 5714 120000 6040 120018
rect -402 119976 -137 119988
rect -402 119936 -390 119976
rect -348 119936 -137 119976
rect -402 119922 -137 119936
rect -589 119909 -499 119915
rect -589 119855 -577 119909
rect -511 119873 -499 119909
rect -511 119855 -241 119873
rect -589 119849 -241 119855
rect -577 119807 -241 119849
rect -963 119670 -336 119680
rect -963 119628 -388 119670
rect -352 119628 -336 119670
rect -963 119614 -336 119628
rect -963 118549 -897 119614
rect -835 119552 -764 119569
rect -835 119516 -820 119552
rect -782 119516 -764 119552
rect -835 119498 -764 119516
rect -532 119534 -438 119540
rect -829 118656 -770 119498
rect -532 119456 -524 119534
rect -446 119456 -438 119534
rect -532 119450 -438 119456
rect -307 119283 -241 119807
rect -545 119277 -241 119283
rect -545 119223 -533 119277
rect -479 119223 -241 119277
rect -545 119217 -241 119223
rect -203 119175 -137 119922
rect 5714 119926 6040 119944
rect 5714 119876 6015 119926
rect 6032 119876 6040 119926
rect 5714 119858 6040 119876
rect 5714 119784 6040 119802
rect 5714 119734 6015 119784
rect 6032 119734 6040 119784
rect 5714 119716 6040 119734
rect 5714 119642 6040 119660
rect 5714 119592 6015 119642
rect 6032 119592 6040 119642
rect 5714 119574 6040 119592
rect 5714 119500 6040 119518
rect 5714 119450 6015 119500
rect 6032 119450 6040 119500
rect 5714 119432 6040 119450
rect 5714 119358 6040 119376
rect 5714 119308 6015 119358
rect 6032 119308 6040 119358
rect 5714 119290 6040 119308
rect -545 119169 -137 119175
rect -545 119115 -533 119169
rect -479 119115 -137 119169
rect 5714 119216 6040 119234
rect 5714 119166 6015 119216
rect 6032 119166 6040 119216
rect 5714 119148 6040 119166
rect -545 119109 -137 119115
rect 5714 119074 6040 119092
rect 5714 119024 6015 119074
rect 6032 119024 6040 119074
rect 5714 119006 6040 119024
rect 5714 118932 6040 118950
rect 5714 118882 6015 118932
rect 6032 118882 6040 118932
rect 5714 118864 6040 118882
rect -637 118827 -571 118833
rect -637 118755 -571 118761
rect 5714 118790 6040 118808
rect 5714 118740 6015 118790
rect 6032 118740 6040 118790
rect 5714 118722 6040 118740
rect -829 118597 -503 118656
rect 5714 118648 6040 118666
rect 5714 118598 6015 118648
rect 6032 118598 6040 118648
rect 5714 118580 6040 118598
rect -963 118483 -701 118549
rect 5714 118506 6040 118524
rect 5714 118456 6015 118506
rect 6032 118456 6040 118506
rect 5714 118438 6040 118456
rect -626 118425 -546 118432
rect -626 118359 -619 118425
rect -553 118359 -546 118425
rect -626 118352 -546 118359
rect 5714 118364 6040 118382
rect 5714 118314 6015 118364
rect 6032 118314 6040 118364
rect 5714 118296 6040 118314
rect 5714 118222 6040 118240
rect -644 118191 -564 118198
rect -644 118125 -637 118191
rect -571 118125 -564 118191
rect 5714 118172 6015 118222
rect 6032 118172 6040 118222
rect 5714 118154 6040 118172
rect -644 118118 -564 118125
rect 5714 118080 6040 118098
rect 5714 118030 6015 118080
rect 6032 118030 6040 118080
rect 5714 118012 6040 118030
rect 5714 117938 6040 117956
rect 5714 117888 6015 117938
rect 6032 117888 6040 117938
rect 5714 117870 6040 117888
rect -634 117811 -538 117818
rect -634 117729 -627 117811
rect -545 117729 -538 117811
rect -634 117722 -538 117729
rect 5714 117796 6040 117814
rect 5714 117746 6015 117796
rect 6032 117746 6040 117796
rect 5714 117728 6040 117746
rect 5714 117654 6040 117672
rect 5714 117604 6015 117654
rect 6032 117604 6040 117654
rect 5714 117586 6040 117604
rect 5714 117512 6040 117530
rect 5714 117462 6015 117512
rect 6032 117462 6040 117512
rect 5714 117444 6040 117462
rect -477 117376 -411 117382
rect -477 117304 -411 117310
rect 5714 117370 6040 117388
rect 5714 117320 6015 117370
rect 6032 117320 6040 117370
rect 5714 117302 6040 117320
rect 5714 117228 6040 117246
rect 5714 117178 6015 117228
rect 6032 117178 6040 117228
rect 5714 117160 6040 117178
rect 5714 117086 6040 117104
rect 5714 117036 6015 117086
rect 6032 117036 6040 117086
rect 5714 117018 6040 117036
rect 5714 116944 6040 116962
rect 5714 116894 6015 116944
rect 6032 116894 6040 116944
rect 5714 116876 6040 116894
rect 5714 116802 6040 116820
rect 5714 116752 6015 116802
rect 6032 116752 6040 116802
rect 5714 116734 6040 116752
rect 5714 116660 6040 116678
rect 5714 116610 6015 116660
rect 6032 116610 6040 116660
rect 5714 116592 6040 116610
rect 5714 116518 6040 116536
rect 5714 116468 6015 116518
rect 6032 116468 6040 116518
rect 5714 116450 6040 116468
rect 5714 116376 6040 116394
rect 5714 116326 6015 116376
rect 6032 116326 6040 116376
rect 5714 116308 6040 116326
rect 5714 116234 6040 116252
rect 5714 116184 6015 116234
rect 6032 116184 6040 116234
rect 5714 116166 6040 116184
rect 5714 116092 6040 116110
rect 5714 116042 6015 116092
rect 6032 116042 6040 116092
rect 5714 116024 6040 116042
rect 5714 115950 6040 115968
rect 5714 115900 6015 115950
rect 6032 115900 6040 115950
rect 5714 115882 6040 115900
rect 5714 115808 6040 115826
rect 5714 115758 6015 115808
rect 6032 115758 6040 115808
rect 5714 115740 6040 115758
rect 5714 115666 6040 115684
rect 5714 115616 6015 115666
rect 6032 115616 6040 115666
rect 5714 115598 6040 115616
rect 5714 115524 6040 115542
rect 5714 115474 6015 115524
rect 6032 115474 6040 115524
rect 5714 115456 6040 115474
rect 5714 115382 6040 115400
rect 5714 115332 6015 115382
rect 6032 115332 6040 115382
rect 5714 115314 6040 115332
rect 5714 115240 6040 115258
rect 5714 115190 6015 115240
rect 6032 115190 6040 115240
rect 5714 115172 6040 115190
rect 5714 115098 6040 115116
rect 5714 115048 6015 115098
rect 6032 115048 6040 115098
rect 5714 115030 6040 115048
rect 5714 114956 6040 114974
rect 5714 114906 6015 114956
rect 6032 114906 6040 114956
rect 5714 114888 6040 114906
rect 5714 114814 6040 114832
rect 5714 114764 6015 114814
rect 6032 114764 6040 114814
rect 5714 114746 6040 114764
rect 5714 114672 6040 114690
rect 5714 114622 6015 114672
rect 6032 114622 6040 114672
rect 5714 114604 6040 114622
rect 5714 114530 6040 114548
rect 5714 114480 6015 114530
rect 6032 114480 6040 114530
rect 5714 114462 6040 114480
rect -412 114390 -346 114400
rect -412 114316 -398 114390
rect 5714 114388 6040 114406
rect -346 114316 -335 114365
rect 5714 114338 6015 114388
rect 6032 114338 6040 114388
rect 5714 114320 6040 114338
rect -401 114299 -335 114316
rect 5714 114246 6040 114264
rect 5714 114196 6015 114246
rect 6032 114196 6040 114246
rect 5714 114178 6040 114196
rect 5714 114104 6040 114122
rect 5714 114054 6015 114104
rect 6032 114054 6040 114104
rect 5714 114036 6040 114054
rect 5714 113962 6040 113980
rect 5714 113912 6015 113962
rect 6032 113912 6040 113962
rect 5714 113894 6040 113912
rect 5714 113820 6040 113838
rect 5714 113770 6015 113820
rect 6032 113770 6040 113820
rect 5714 113752 6040 113770
rect 5714 113678 6040 113696
rect 5714 113628 6015 113678
rect 6032 113628 6040 113678
rect 5714 113610 6040 113628
rect 5714 113536 6040 113554
rect 5714 113486 6015 113536
rect 6032 113486 6040 113536
rect 5714 113468 6040 113486
rect 5714 113394 6040 113412
rect 5714 113344 6015 113394
rect 6032 113344 6040 113394
rect 5714 113326 6040 113344
rect 5714 113252 6040 113270
rect 5714 113202 6015 113252
rect 6032 113202 6040 113252
rect 5714 113184 6040 113202
rect 5714 113110 6040 113128
rect 5714 113060 6015 113110
rect 6032 113060 6040 113110
rect 5714 113042 6040 113060
rect 5714 112968 6040 112986
rect 5714 112918 6015 112968
rect 6032 112918 6040 112968
rect 5714 112900 6040 112918
rect 5714 112826 6040 112844
rect 5714 112776 6015 112826
rect 6032 112776 6040 112826
rect 5714 112758 6040 112776
rect 5714 112684 6040 112702
rect 5714 112634 6015 112684
rect 6032 112634 6040 112684
rect 5714 112616 6040 112634
rect 5714 112542 6040 112560
rect 5714 112492 6015 112542
rect 6032 112492 6040 112542
rect 5714 112474 6040 112492
rect 5714 112400 6040 112418
rect 5714 112350 6015 112400
rect 6032 112350 6040 112400
rect 5714 112332 6040 112350
rect 5714 112258 6040 112276
rect 5714 112208 6015 112258
rect 6032 112208 6040 112258
rect 5714 112190 6040 112208
rect 5714 112116 6040 112134
rect 5714 112066 6015 112116
rect 6032 112066 6040 112116
rect 5714 112048 6040 112066
rect 5714 111974 6040 111992
rect 5714 111924 6015 111974
rect 6032 111924 6040 111974
rect 5714 111906 6040 111924
rect 5714 111832 6040 111850
rect 5714 111782 6015 111832
rect 6032 111782 6040 111832
rect 5714 111764 6040 111782
rect 5714 111690 6040 111708
rect 5714 111640 6015 111690
rect 6032 111640 6040 111690
rect 5714 111622 6040 111640
rect 5714 111548 6040 111566
rect 5714 111498 6015 111548
rect 6032 111498 6040 111548
rect 5714 111480 6040 111498
rect 5714 111406 6040 111424
rect 5714 111356 6015 111406
rect 6032 111356 6040 111406
rect 5714 111338 6040 111356
rect 5714 111264 6040 111282
rect 5714 111214 6015 111264
rect 6032 111214 6040 111264
rect 5714 111196 6040 111214
rect 5714 111122 6040 111140
rect 5714 111072 6015 111122
rect 6032 111072 6040 111122
rect 5714 111054 6040 111072
rect 5714 110980 6040 110998
rect 5714 110930 6015 110980
rect 6032 110930 6040 110980
rect 5714 110912 6040 110930
rect 5714 110838 6040 110856
rect 5714 110788 6015 110838
rect 6032 110788 6040 110838
rect 5714 110770 6040 110788
rect 5714 110696 6040 110714
rect 5714 110646 6015 110696
rect 6032 110646 6040 110696
rect 5714 110628 6040 110646
rect 5714 110554 6040 110572
rect 5714 110504 6015 110554
rect 6032 110504 6040 110554
rect 5714 110486 6040 110504
rect 5714 110412 6040 110430
rect 5714 110362 6015 110412
rect 6032 110362 6040 110412
rect 5714 110344 6040 110362
rect 5714 110270 6040 110288
rect 5714 110220 6015 110270
rect 6032 110220 6040 110270
rect 5714 110202 6040 110220
rect 5714 110128 6040 110146
rect 5714 110078 6015 110128
rect 6032 110078 6040 110128
rect 5714 110060 6040 110078
rect 5714 109986 6040 110004
rect 5714 109936 6015 109986
rect 6032 109936 6040 109986
rect 5714 109918 6040 109936
rect 5714 109844 6040 109862
rect 5714 109794 6015 109844
rect 6032 109794 6040 109844
rect 5714 109776 6040 109794
rect 5714 109702 6040 109720
rect 5714 109652 6015 109702
rect 6032 109652 6040 109702
rect 5714 109634 6040 109652
rect 5714 109560 6040 109578
rect 5714 109510 6015 109560
rect 6032 109510 6040 109560
rect 5714 109492 6040 109510
rect 5714 109418 6040 109436
rect 5714 109368 6015 109418
rect 6032 109368 6040 109418
rect 5714 109350 6040 109368
rect 5714 109276 6040 109294
rect 5714 109226 6015 109276
rect 6032 109226 6040 109276
rect 5714 109208 6040 109226
rect 5714 109134 6040 109152
rect 5714 109084 6015 109134
rect 6032 109084 6040 109134
rect 5714 109066 6040 109084
rect 5714 108992 6040 109010
rect 5714 108942 6015 108992
rect 6032 108942 6040 108992
rect 5714 108924 6040 108942
rect 5714 108850 6040 108868
rect 5714 108800 6015 108850
rect 6032 108800 6040 108850
rect 5714 108782 6040 108800
rect 5714 108708 6040 108726
rect 5714 108658 6015 108708
rect 6032 108658 6040 108708
rect 5714 108640 6040 108658
rect 5714 108566 6040 108584
rect 5714 108516 6015 108566
rect 6032 108516 6040 108566
rect 5714 108498 6040 108516
rect 5714 108424 6040 108442
rect 5714 108374 6015 108424
rect 6032 108374 6040 108424
rect 5714 108356 6040 108374
rect 5714 108282 6040 108300
rect 5714 108232 6015 108282
rect 6032 108232 6040 108282
rect 5714 108214 6040 108232
rect 5714 108140 6040 108158
rect 5714 108090 6015 108140
rect 6032 108090 6040 108140
rect 5714 108072 6040 108090
rect 5714 107998 6040 108016
rect 5714 107948 6015 107998
rect 6032 107948 6040 107998
rect 5714 107930 6040 107948
rect -406 107894 -332 107904
rect -406 107814 -394 107894
rect -338 107814 -332 107894
rect -406 107802 -332 107814
rect 5714 107856 6040 107874
rect 5714 107806 6015 107856
rect 6032 107806 6040 107856
rect 5714 107788 6040 107806
rect 5714 107714 6040 107732
rect 5714 107664 6015 107714
rect 6032 107664 6040 107714
rect 5714 107646 6040 107664
rect 5714 107572 6040 107590
rect 5714 107522 6015 107572
rect 6032 107522 6040 107572
rect 5714 107504 6040 107522
rect 5714 107430 6040 107448
rect 5714 107380 6015 107430
rect 6032 107380 6040 107430
rect 5714 107362 6040 107380
rect 5714 107288 6040 107306
rect 5714 107238 6015 107288
rect 6032 107238 6040 107288
rect 5714 107220 6040 107238
rect 5714 107146 6040 107164
rect 5714 107096 6015 107146
rect 6032 107096 6040 107146
rect 5714 107078 6040 107096
rect 5714 107004 6040 107022
rect 5714 106954 6015 107004
rect 6032 106954 6040 107004
rect 5714 106936 6040 106954
rect 5714 106862 6040 106880
rect 5714 106812 6015 106862
rect 6032 106812 6040 106862
rect 5714 106794 6040 106812
rect 5714 106720 6040 106738
rect 5714 106670 6015 106720
rect 6032 106670 6040 106720
rect 5714 106652 6040 106670
rect 5714 106578 6040 106596
rect 5714 106528 6015 106578
rect 6032 106528 6040 106578
rect 5714 106510 6040 106528
rect 5714 106436 6040 106454
rect 5714 106386 6015 106436
rect 6032 106386 6040 106436
rect 5714 106368 6040 106386
rect 5714 106294 6040 106312
rect 5714 106244 6015 106294
rect 6032 106244 6040 106294
rect 5714 106226 6040 106244
rect 5714 106152 6040 106170
rect 5714 106102 6015 106152
rect 6032 106102 6040 106152
rect 5714 106084 6040 106102
rect 5714 106010 6040 106028
rect 5714 105960 6015 106010
rect 6032 105960 6040 106010
rect 5714 105942 6040 105960
rect 5714 105868 6040 105886
rect 5714 105818 6015 105868
rect 6032 105818 6040 105868
rect 5714 105800 6040 105818
rect 5714 105726 6040 105744
rect 5714 105676 6015 105726
rect 6032 105676 6040 105726
rect 5714 105658 6040 105676
rect 5714 105584 6040 105602
rect 5714 105534 6015 105584
rect 6032 105534 6040 105584
rect 5714 105516 6040 105534
rect 5714 105442 6040 105460
rect 5714 105392 6015 105442
rect 6032 105392 6040 105442
rect 5714 105374 6040 105392
rect 5714 105300 6040 105318
rect 5714 105250 6015 105300
rect 6032 105250 6040 105300
rect 5714 105232 6040 105250
rect 5714 105158 6040 105176
rect 5714 105108 6015 105158
rect 6032 105108 6040 105158
rect 5714 105090 6040 105108
rect 5714 105016 6040 105034
rect 5714 104966 6015 105016
rect 6032 104966 6040 105016
rect 5714 104948 6040 104966
rect 5714 104874 6040 104892
rect 5714 104824 6015 104874
rect 6032 104824 6040 104874
rect 5714 104806 6040 104824
rect 5714 104732 6040 104750
rect 5714 104682 6015 104732
rect 6032 104682 6040 104732
rect 5714 104664 6040 104682
rect 5714 104590 6040 104608
rect 5714 104540 6015 104590
rect 6032 104540 6040 104590
rect 5714 104522 6040 104540
rect 5714 104448 6040 104466
rect 5714 104398 6015 104448
rect 6032 104398 6040 104448
rect 5714 104380 6040 104398
rect 5714 104306 6040 104324
rect 5714 104256 6015 104306
rect 6032 104256 6040 104306
rect 5714 104238 6040 104256
rect 5714 104164 6040 104182
rect 5714 104114 6015 104164
rect 6032 104114 6040 104164
rect 5714 104096 6040 104114
rect 5714 104022 6040 104040
rect 5714 103972 6015 104022
rect 6032 103972 6040 104022
rect 5714 103954 6040 103972
rect 5714 103880 6040 103898
rect 5714 103830 6015 103880
rect 6032 103830 6040 103880
rect 5714 103812 6040 103830
rect 5714 103738 6040 103756
rect 5714 103688 6015 103738
rect 6032 103688 6040 103738
rect 5714 103670 6040 103688
rect 5714 103596 6040 103614
rect 5714 103546 6015 103596
rect 6032 103546 6040 103596
rect 5714 103528 6040 103546
rect 5714 103454 6040 103472
rect 5714 103404 6015 103454
rect 6032 103404 6040 103454
rect 5714 103386 6040 103404
rect 5714 103312 6040 103330
rect 5714 103262 6015 103312
rect 6032 103262 6040 103312
rect 5714 103244 6040 103262
rect 5714 103170 6040 103188
rect 5714 103120 6015 103170
rect 6032 103120 6040 103170
rect 5714 103102 6040 103120
rect 5714 103028 6040 103046
rect 5714 102978 6015 103028
rect 6032 102978 6040 103028
rect 5714 102960 6040 102978
rect 5714 102886 6040 102904
rect 5714 102836 6015 102886
rect 6032 102836 6040 102886
rect 5714 102818 6040 102836
rect 5714 102744 6040 102762
rect 5714 102694 6015 102744
rect 6032 102694 6040 102744
rect 5714 102676 6040 102694
rect 5714 102602 6040 102620
rect 5714 102552 6015 102602
rect 6032 102552 6040 102602
rect 5714 102534 6040 102552
rect 5714 102460 6040 102478
rect 5714 102410 6015 102460
rect 6032 102410 6040 102460
rect 5714 102392 6040 102410
rect 5714 102318 6040 102336
rect 5714 102268 6015 102318
rect 6032 102268 6040 102318
rect 5714 102250 6040 102268
rect 5714 102176 6040 102194
rect 5714 102126 6015 102176
rect 6032 102126 6040 102176
rect 5714 102108 6040 102126
rect 5714 102034 6040 102052
rect 5714 101984 6015 102034
rect 6032 101984 6040 102034
rect 5714 101966 6040 101984
rect 5714 101892 6040 101910
rect 5714 101842 6015 101892
rect 6032 101842 6040 101892
rect 5714 101824 6040 101842
rect 5714 101750 6040 101768
rect 5714 101700 6015 101750
rect 6032 101700 6040 101750
rect 5714 101682 6040 101700
rect 5714 101608 6040 101626
rect 5714 101558 6015 101608
rect 6032 101558 6040 101608
rect 5714 101540 6040 101558
rect 5714 101466 6040 101484
rect 5714 101416 6015 101466
rect 6032 101416 6040 101466
rect 5714 101398 6040 101416
rect 5714 101324 6040 101342
rect 5714 101274 6015 101324
rect 6032 101274 6040 101324
rect 5714 101256 6040 101274
rect 5714 101182 6040 101200
rect 5714 101132 6015 101182
rect 6032 101132 6040 101182
rect 5714 101114 6040 101132
rect 5714 101040 6040 101058
rect 5714 100990 6015 101040
rect 6032 100990 6040 101040
rect 5714 100972 6040 100990
rect 5714 100898 6040 100916
rect 5714 100848 6015 100898
rect 6032 100848 6040 100898
rect 5714 100830 6040 100848
rect 5714 100756 6040 100774
rect 5714 100706 6015 100756
rect 6032 100706 6040 100756
rect 5714 100688 6040 100706
rect 5714 100614 6040 100632
rect 5714 100564 6015 100614
rect 6032 100564 6040 100614
rect 5714 100546 6040 100564
rect 5714 100472 6040 100490
rect 5714 100422 6015 100472
rect 6032 100422 6040 100472
rect 5714 100404 6040 100422
rect 5714 100330 6040 100348
rect 5714 100280 6015 100330
rect 6032 100280 6040 100330
rect 5714 100262 6040 100280
rect 5714 100188 6040 100206
rect 5714 100138 6015 100188
rect 6032 100138 6040 100188
rect 5714 100120 6040 100138
rect 5714 100046 6040 100064
rect 5714 99996 6015 100046
rect 6032 99996 6040 100046
rect 5714 99978 6040 99996
rect 5714 99904 6040 99922
rect 5714 99854 6015 99904
rect 6032 99854 6040 99904
rect 5714 99836 6040 99854
rect 5714 99762 6040 99780
rect 5714 99712 6015 99762
rect 6032 99712 6040 99762
rect 5714 99694 6040 99712
rect 5714 99620 6040 99638
rect 5714 99570 6015 99620
rect 6032 99570 6040 99620
rect 5714 99552 6040 99570
rect 5714 99478 6040 99496
rect 5714 99428 6015 99478
rect 6032 99428 6040 99478
rect 5714 99410 6040 99428
rect 5714 99336 6040 99354
rect 5714 99286 6015 99336
rect 6032 99286 6040 99336
rect 5714 99268 6040 99286
rect 5714 99194 6040 99212
rect 5714 99144 6015 99194
rect 6032 99144 6040 99194
rect 5714 99126 6040 99144
rect 5714 99052 6040 99070
rect 5714 99002 6015 99052
rect 6032 99002 6040 99052
rect 5714 98984 6040 99002
rect 5714 98910 6040 98928
rect 5714 98860 6015 98910
rect 6032 98860 6040 98910
rect 5714 98842 6040 98860
rect 5714 98768 6040 98786
rect 5714 98718 6015 98768
rect 6032 98718 6040 98768
rect 5714 98700 6040 98718
rect 5714 98626 6040 98644
rect 5714 98576 6015 98626
rect 6032 98576 6040 98626
rect 5714 98558 6040 98576
rect 5714 98484 6040 98502
rect 5714 98434 6015 98484
rect 6032 98434 6040 98484
rect 5714 98416 6040 98434
rect 5714 98342 6040 98360
rect 5714 98292 6015 98342
rect 6032 98292 6040 98342
rect 5714 98274 6040 98292
rect 5714 98200 6040 98218
rect 5714 98150 6015 98200
rect 6032 98150 6040 98200
rect 5714 98132 6040 98150
rect 5714 98058 6040 98076
rect 5714 98008 6015 98058
rect 6032 98008 6040 98058
rect 5714 97990 6040 98008
rect 5714 97916 6040 97934
rect 5714 97866 6015 97916
rect 6032 97866 6040 97916
rect 5714 97848 6040 97866
rect 5714 97774 6040 97792
rect 5714 97724 6015 97774
rect 6032 97724 6040 97774
rect 5714 97706 6040 97724
rect 5714 97632 6040 97650
rect 5714 97582 6015 97632
rect 6032 97582 6040 97632
rect 5714 97564 6040 97582
rect 5714 97490 6040 97508
rect 5714 97440 6015 97490
rect 6032 97440 6040 97490
rect 5714 97422 6040 97440
rect 5714 97348 6040 97366
rect 5714 97298 6015 97348
rect 6032 97298 6040 97348
rect 5714 97280 6040 97298
rect 5714 97206 6040 97224
rect 5714 97156 6015 97206
rect 6032 97156 6040 97206
rect 5714 97138 6040 97156
rect 5714 97064 6040 97082
rect 5714 97014 6015 97064
rect 6032 97014 6040 97064
rect 5714 96996 6040 97014
rect 5714 96922 6040 96940
rect 5714 96872 6015 96922
rect 6032 96872 6040 96922
rect 5714 96854 6040 96872
rect 5714 96780 6040 96798
rect 5714 96730 6015 96780
rect 6032 96730 6040 96780
rect 5714 96712 6040 96730
rect 5714 96638 6040 96656
rect 5714 96588 6015 96638
rect 6032 96588 6040 96638
rect 5714 96570 6040 96588
rect 5714 96496 6040 96514
rect 5714 96446 6015 96496
rect 6032 96446 6040 96496
rect 5714 96428 6040 96446
rect 5714 96354 6040 96372
rect 5714 96304 6015 96354
rect 6032 96304 6040 96354
rect 5714 96286 6040 96304
rect 5714 96212 6040 96230
rect 5714 96162 6015 96212
rect 6032 96162 6040 96212
rect 5714 96144 6040 96162
rect 5714 96070 6040 96088
rect 5714 96020 6015 96070
rect 6032 96020 6040 96070
rect 5714 96002 6040 96020
rect 5714 95928 6040 95946
rect 5714 95878 6015 95928
rect 6032 95878 6040 95928
rect 5714 95860 6040 95878
rect 5714 95786 6040 95804
rect 5714 95736 6015 95786
rect 6032 95736 6040 95786
rect 5714 95718 6040 95736
rect 5714 95644 6040 95662
rect 5714 95594 6015 95644
rect 6032 95594 6040 95644
rect 5714 95576 6040 95594
rect 5714 95502 6040 95520
rect 5714 95452 6015 95502
rect 6032 95452 6040 95502
rect 5714 95434 6040 95452
rect 5714 95360 6040 95378
rect 5714 95310 6015 95360
rect 6032 95310 6040 95360
rect 5714 95292 6040 95310
rect 5714 95218 6040 95236
rect 5714 95168 6015 95218
rect 6032 95168 6040 95218
rect 5714 95150 6040 95168
rect 5714 95076 6040 95094
rect 5714 95026 6015 95076
rect 6032 95026 6040 95076
rect 5714 95008 6040 95026
rect 5714 94934 6040 94952
rect 5714 94884 6015 94934
rect 6032 94884 6040 94934
rect 5714 94866 6040 94884
rect 5714 94792 6040 94810
rect 5714 94742 6015 94792
rect 6032 94742 6040 94792
rect 5714 94724 6040 94742
rect 5714 94650 6040 94668
rect 5714 94600 6015 94650
rect 6032 94600 6040 94650
rect 5714 94582 6040 94600
rect 5714 94508 6040 94526
rect 5714 94458 6015 94508
rect 6032 94458 6040 94508
rect 5714 94440 6040 94458
rect 5714 94366 6040 94384
rect 5714 94316 6015 94366
rect 6032 94316 6040 94366
rect 5714 94298 6040 94316
rect 5714 94224 6040 94242
rect 5714 94174 6015 94224
rect 6032 94174 6040 94224
rect 5714 94156 6040 94174
rect 5714 94082 6040 94100
rect 5714 94032 6015 94082
rect 6032 94032 6040 94082
rect 5714 94014 6040 94032
rect 5714 93940 6040 93958
rect 5714 93890 6015 93940
rect 6032 93890 6040 93940
rect 5714 93872 6040 93890
rect 5714 93798 6040 93816
rect 5714 93748 6015 93798
rect 6032 93748 6040 93798
rect 5714 93730 6040 93748
rect 5714 93656 6040 93674
rect 5714 93606 6015 93656
rect 6032 93606 6040 93656
rect 5714 93588 6040 93606
rect 5714 93514 6040 93532
rect 5714 93464 6015 93514
rect 6032 93464 6040 93514
rect 5714 93446 6040 93464
rect 5714 93372 6040 93390
rect 5714 93322 6015 93372
rect 6032 93322 6040 93372
rect 5714 93304 6040 93322
rect 5714 93230 6040 93248
rect 5714 93180 6015 93230
rect 6032 93180 6040 93230
rect 5714 93162 6040 93180
rect 5714 93088 6040 93106
rect 5714 93038 6015 93088
rect 6032 93038 6040 93088
rect 5714 93020 6040 93038
rect 5714 92946 6040 92964
rect 5714 92896 6015 92946
rect 6032 92896 6040 92946
rect 5714 92878 6040 92896
rect 5714 92804 6040 92822
rect 5714 92754 6015 92804
rect 6032 92754 6040 92804
rect 5714 92736 6040 92754
rect 5714 92662 6040 92680
rect 5714 92612 6015 92662
rect 6032 92612 6040 92662
rect 5714 92594 6040 92612
rect 5714 92520 6040 92538
rect 5714 92470 6015 92520
rect 6032 92470 6040 92520
rect 5714 92452 6040 92470
rect 5714 92378 6040 92396
rect 5714 92328 6015 92378
rect 6032 92328 6040 92378
rect 5714 92310 6040 92328
rect 5714 92236 6040 92254
rect 5714 92186 6015 92236
rect 6032 92186 6040 92236
rect 5714 92168 6040 92186
rect 5714 92094 6040 92112
rect 5714 92044 6015 92094
rect 6032 92044 6040 92094
rect 5714 92026 6040 92044
rect 5714 91952 6040 91970
rect 5714 91902 6015 91952
rect 6032 91902 6040 91952
rect 5714 91884 6040 91902
rect 5714 91810 6040 91828
rect 5714 91760 6015 91810
rect 6032 91760 6040 91810
rect 5714 91742 6040 91760
rect 5714 91668 6040 91686
rect 5714 91618 6015 91668
rect 6032 91618 6040 91668
rect 5714 91600 6040 91618
rect 5714 91526 6040 91544
rect 5714 91476 6015 91526
rect 6032 91476 6040 91526
rect 5714 91458 6040 91476
rect 5714 91384 6040 91402
rect 5714 91334 6015 91384
rect 6032 91334 6040 91384
rect 5714 91316 6040 91334
rect 5714 91242 6040 91260
rect 5714 91192 6015 91242
rect 6032 91192 6040 91242
rect 5714 91174 6040 91192
rect 5714 91100 6040 91118
rect 5714 91050 6015 91100
rect 6032 91050 6040 91100
rect 5714 91032 6040 91050
rect 5714 90958 6040 90976
rect 5714 90908 6015 90958
rect 6032 90908 6040 90958
rect 5714 90890 6040 90908
rect 5714 90816 6040 90834
rect 5714 90766 6015 90816
rect 6032 90766 6040 90816
rect 5714 90748 6040 90766
rect 5714 90674 6040 90692
rect 5714 90624 6015 90674
rect 6032 90624 6040 90674
rect 5714 90606 6040 90624
rect 5714 90532 6040 90550
rect 5714 90482 6015 90532
rect 6032 90482 6040 90532
rect 5714 90464 6040 90482
rect 5714 90390 6040 90408
rect 5714 90340 6015 90390
rect 6032 90340 6040 90390
rect 5714 90322 6040 90340
rect 5714 90248 6040 90266
rect 5714 90198 6015 90248
rect 6032 90198 6040 90248
rect 5714 90180 6040 90198
rect 5714 90106 6040 90124
rect 5714 90056 6015 90106
rect 6032 90056 6040 90106
rect 5714 90038 6040 90056
rect 5714 89964 6040 89982
rect 5714 89914 6015 89964
rect 6032 89914 6040 89964
rect 5714 89896 6040 89914
rect 5714 89822 6040 89840
rect 5714 89772 6015 89822
rect 6032 89772 6040 89822
rect 5714 89754 6040 89772
rect 5714 89680 6040 89698
rect 5714 89630 6015 89680
rect 6032 89630 6040 89680
rect 5714 89612 6040 89630
rect 5714 89538 6040 89556
rect 5714 89488 6015 89538
rect 6032 89488 6040 89538
rect 5714 89470 6040 89488
rect 5714 89396 6040 89414
rect 5714 89346 6015 89396
rect 6032 89346 6040 89396
rect 5714 89328 6040 89346
rect 5714 89254 6040 89272
rect 5714 89204 6015 89254
rect 6032 89204 6040 89254
rect 5714 89186 6040 89204
rect 5714 89112 6040 89130
rect 5714 89062 6015 89112
rect 6032 89062 6040 89112
rect 5714 89044 6040 89062
rect 5714 88970 6040 88988
rect 5714 88920 6015 88970
rect 6032 88920 6040 88970
rect 5714 88902 6040 88920
rect 5714 88828 6040 88846
rect 5714 88778 6015 88828
rect 6032 88778 6040 88828
rect 5714 88760 6040 88778
rect 5714 88686 6040 88704
rect 5714 88636 6015 88686
rect 6032 88636 6040 88686
rect 5714 88618 6040 88636
rect 5714 88544 6040 88562
rect 5714 88494 6015 88544
rect 6032 88494 6040 88544
rect 5714 88476 6040 88494
rect 5714 88402 6040 88420
rect 5714 88352 6015 88402
rect 6032 88352 6040 88402
rect 5714 88334 6040 88352
rect 5714 88260 6040 88278
rect 5714 88210 6015 88260
rect 6032 88210 6040 88260
rect 5714 88192 6040 88210
rect 5714 88118 6040 88136
rect 5714 88068 6015 88118
rect 6032 88068 6040 88118
rect 5714 88050 6040 88068
rect 5714 87976 6040 87994
rect 5714 87926 6015 87976
rect 6032 87926 6040 87976
rect 5714 87908 6040 87926
rect 5714 87834 6040 87852
rect 5714 87784 6015 87834
rect 6032 87784 6040 87834
rect 5714 87766 6040 87784
rect 5714 87692 6040 87710
rect 5714 87642 6015 87692
rect 6032 87642 6040 87692
rect 5714 87624 6040 87642
rect 5714 87550 6040 87568
rect 5714 87500 6015 87550
rect 6032 87500 6040 87550
rect 5714 87482 6040 87500
rect 5714 87408 6040 87426
rect 5714 87358 6015 87408
rect 6032 87358 6040 87408
rect 5714 87340 6040 87358
rect 5714 87266 6040 87284
rect 5714 87216 6015 87266
rect 6032 87216 6040 87266
rect 5714 87198 6040 87216
rect 5714 87124 6040 87142
rect 5714 87074 6015 87124
rect 6032 87074 6040 87124
rect 5714 87056 6040 87074
rect 5714 86982 6040 87000
rect 5714 86932 6015 86982
rect 6032 86932 6040 86982
rect 5714 86914 6040 86932
rect 5714 86840 6040 86858
rect 5714 86790 6015 86840
rect 6032 86790 6040 86840
rect 5714 86772 6040 86790
rect 5714 86698 6040 86716
rect 5714 86648 6015 86698
rect 6032 86648 6040 86698
rect 5714 86630 6040 86648
rect 5714 86556 6040 86574
rect 5714 86506 6015 86556
rect 6032 86506 6040 86556
rect 5714 86488 6040 86506
rect 5714 86414 6040 86432
rect 5714 86364 6015 86414
rect 6032 86364 6040 86414
rect 5714 86346 6040 86364
rect 5714 86272 6040 86290
rect 5714 86222 6015 86272
rect 6032 86222 6040 86272
rect 5714 86204 6040 86222
rect 5714 86130 6040 86148
rect 5714 86080 6015 86130
rect 6032 86080 6040 86130
rect 5714 86062 6040 86080
rect 5714 85988 6040 86006
rect 5714 85938 6015 85988
rect 6032 85938 6040 85988
rect 5714 85920 6040 85938
rect 5714 85846 6040 85864
rect 5714 85796 6015 85846
rect 6032 85796 6040 85846
rect 5714 85778 6040 85796
rect 5714 85704 6040 85722
rect 5714 85654 6015 85704
rect 6032 85654 6040 85704
rect 5714 85636 6040 85654
rect 5714 85562 6040 85580
rect 5714 85512 6015 85562
rect 6032 85512 6040 85562
rect 5714 85494 6040 85512
rect 5714 85420 6040 85438
rect 5714 85370 6015 85420
rect 6032 85370 6040 85420
rect 5714 85352 6040 85370
rect 5714 85278 6040 85296
rect 5714 85228 6015 85278
rect 6032 85228 6040 85278
rect 5714 85210 6040 85228
rect 5714 85136 6040 85154
rect 5714 85086 6015 85136
rect 6032 85086 6040 85136
rect 5714 85068 6040 85086
rect 5714 84994 6040 85012
rect 5714 84944 6015 84994
rect 6032 84944 6040 84994
rect 5714 84926 6040 84944
rect 5714 84852 6040 84870
rect 5714 84802 6015 84852
rect 6032 84802 6040 84852
rect 5714 84784 6040 84802
rect 5714 84710 6040 84728
rect 5714 84660 6015 84710
rect 6032 84660 6040 84710
rect 5714 84642 6040 84660
rect 5714 84568 6040 84586
rect 5714 84518 6015 84568
rect 6032 84518 6040 84568
rect 5714 84500 6040 84518
rect 5714 84426 6040 84444
rect 5714 84376 6015 84426
rect 6032 84376 6040 84426
rect 5714 84358 6040 84376
rect 5714 84284 6040 84302
rect 5714 84234 6015 84284
rect 6032 84234 6040 84284
rect 5714 84216 6040 84234
rect 5714 84142 6040 84160
rect 5714 84092 6015 84142
rect 6032 84092 6040 84142
rect 5714 84074 6040 84092
rect 5714 84000 6040 84018
rect 5714 83950 6015 84000
rect 6032 83950 6040 84000
rect 5714 83932 6040 83950
rect 5714 83858 6040 83876
rect 5714 83808 6015 83858
rect 6032 83808 6040 83858
rect 5714 83790 6040 83808
rect 5714 83716 6040 83734
rect 5714 83666 6015 83716
rect 6032 83666 6040 83716
rect 5714 83648 6040 83666
rect 5714 83574 6040 83592
rect 5714 83524 6015 83574
rect 6032 83524 6040 83574
rect 5714 83506 6040 83524
rect 5714 83432 6040 83450
rect 5714 83382 6015 83432
rect 6032 83382 6040 83432
rect 5714 83364 6040 83382
rect 5714 83290 6040 83308
rect 5714 83240 6015 83290
rect 6032 83240 6040 83290
rect 5714 83222 6040 83240
rect 5714 83148 6040 83166
rect 5714 83098 6015 83148
rect 6032 83098 6040 83148
rect 5714 83080 6040 83098
rect 5714 83006 6040 83024
rect 5714 82956 6015 83006
rect 6032 82956 6040 83006
rect 5714 82938 6040 82956
rect 5714 82864 6040 82882
rect 5714 82814 6015 82864
rect 6032 82814 6040 82864
rect 5714 82796 6040 82814
rect 5714 82722 6040 82740
rect 5714 82672 6015 82722
rect 6032 82672 6040 82722
rect 5714 82654 6040 82672
rect 5714 82580 6040 82598
rect 5714 82530 6015 82580
rect 6032 82530 6040 82580
rect 5714 82512 6040 82530
rect 5714 82438 6040 82456
rect 5714 82388 6015 82438
rect 6032 82388 6040 82438
rect 5714 82370 6040 82388
rect 5714 82296 6040 82314
rect 5714 82246 6015 82296
rect 6032 82246 6040 82296
rect 5714 82228 6040 82246
rect 5714 82154 6040 82172
rect 5714 82104 6015 82154
rect 6032 82104 6040 82154
rect 5714 82086 6040 82104
rect 5714 82012 6040 82030
rect 5714 81962 6015 82012
rect 6032 81962 6040 82012
rect 5714 81944 6040 81962
rect 5714 81870 6040 81888
rect 5714 81820 6015 81870
rect 6032 81820 6040 81870
rect 5714 81802 6040 81820
rect 5714 81728 6040 81746
rect 5714 81678 6015 81728
rect 6032 81678 6040 81728
rect 5714 81660 6040 81678
rect 5714 81586 6040 81604
rect 5714 81536 6015 81586
rect 6032 81536 6040 81586
rect 5714 81518 6040 81536
rect 5714 81444 6040 81462
rect 5714 81394 6015 81444
rect 6032 81394 6040 81444
rect 5714 81376 6040 81394
rect 5714 81302 6040 81320
rect 5714 81252 6015 81302
rect 6032 81252 6040 81302
rect 5714 81234 6040 81252
rect 5714 81160 6040 81178
rect 5714 81110 6015 81160
rect 6032 81110 6040 81160
rect 5714 81092 6040 81110
rect 5714 81018 6040 81036
rect 5714 80968 6015 81018
rect 6032 80968 6040 81018
rect 5714 80950 6040 80968
rect 5714 80876 6040 80894
rect 5714 80826 6015 80876
rect 6032 80826 6040 80876
rect 5714 80808 6040 80826
rect 5714 80734 6040 80752
rect 5714 80684 6015 80734
rect 6032 80684 6040 80734
rect 5714 80666 6040 80684
rect 5714 80592 6040 80610
rect 5714 80542 6015 80592
rect 6032 80542 6040 80592
rect 5714 80524 6040 80542
rect 5714 80450 6040 80468
rect 5714 80400 6015 80450
rect 6032 80400 6040 80450
rect 5714 80382 6040 80400
rect 5714 80308 6040 80326
rect 5714 80258 6015 80308
rect 6032 80258 6040 80308
rect 5714 80240 6040 80258
rect 5714 80166 6040 80184
rect 5714 80116 6015 80166
rect 6032 80116 6040 80166
rect 5714 80098 6040 80116
rect 5714 80024 6040 80042
rect 5714 79974 6015 80024
rect 6032 79974 6040 80024
rect 5714 79956 6040 79974
rect 5714 79882 6040 79900
rect 5714 79832 6015 79882
rect 6032 79832 6040 79882
rect 5714 79814 6040 79832
rect 5714 79740 6040 79758
rect 5714 79690 6015 79740
rect 6032 79690 6040 79740
rect 5714 79672 6040 79690
rect 5714 79598 6040 79616
rect 5714 79548 6015 79598
rect 6032 79548 6040 79598
rect 5714 79530 6040 79548
rect 5714 79456 6040 79474
rect 5714 79406 6015 79456
rect 6032 79406 6040 79456
rect 5714 79388 6040 79406
rect 5714 79314 6040 79332
rect 5714 79264 6015 79314
rect 6032 79264 6040 79314
rect 5714 79246 6040 79264
rect 5714 79172 6040 79190
rect 5714 79122 6015 79172
rect 6032 79122 6040 79172
rect 5714 79104 6040 79122
rect 5714 79030 6040 79048
rect 5714 78980 6015 79030
rect 6032 78980 6040 79030
rect 5714 78962 6040 78980
rect 5714 78888 6040 78906
rect 5714 78838 6015 78888
rect 6032 78838 6040 78888
rect 5714 78820 6040 78838
rect 5714 78746 6040 78764
rect 5714 78696 6015 78746
rect 6032 78696 6040 78746
rect 5714 78678 6040 78696
rect 5714 78604 6040 78622
rect 5714 78554 6015 78604
rect 6032 78554 6040 78604
rect 5714 78536 6040 78554
rect 5714 78462 6040 78480
rect 5714 78412 6015 78462
rect 6032 78412 6040 78462
rect 5714 78394 6040 78412
rect 5714 78320 6040 78338
rect 5714 78270 6015 78320
rect 6032 78270 6040 78320
rect 5714 78252 6040 78270
rect 5714 78178 6040 78196
rect 5714 78128 6015 78178
rect 6032 78128 6040 78178
rect 5714 78110 6040 78128
rect 5714 78036 6040 78054
rect 5714 77986 6015 78036
rect 6032 77986 6040 78036
rect 5714 77968 6040 77986
rect 5714 77894 6040 77912
rect 5714 77844 6015 77894
rect 6032 77844 6040 77894
rect 5714 77826 6040 77844
rect 5714 77752 6040 77770
rect 5714 77702 6015 77752
rect 6032 77702 6040 77752
rect 5714 77684 6040 77702
rect 5714 77610 6040 77628
rect 5714 77560 6015 77610
rect 6032 77560 6040 77610
rect 5714 77542 6040 77560
rect 5714 77468 6040 77486
rect 5714 77418 6015 77468
rect 6032 77418 6040 77468
rect 5714 77400 6040 77418
rect 5714 77326 6040 77344
rect 5714 77276 6015 77326
rect 6032 77276 6040 77326
rect 5714 77258 6040 77276
rect 5714 77184 6040 77202
rect 5714 77134 6015 77184
rect 6032 77134 6040 77184
rect 5714 77116 6040 77134
rect 5714 77042 6040 77060
rect 5714 76992 6015 77042
rect 6032 76992 6040 77042
rect 5714 76974 6040 76992
rect 5714 76900 6040 76918
rect 5714 76850 6015 76900
rect 6032 76850 6040 76900
rect 5714 76832 6040 76850
rect 5714 76758 6040 76776
rect 5714 76708 6015 76758
rect 6032 76708 6040 76758
rect 5714 76690 6040 76708
rect 5714 76616 6040 76634
rect 5714 76566 6015 76616
rect 6032 76566 6040 76616
rect 5714 76548 6040 76566
rect 5714 76474 6040 76492
rect 5714 76424 6015 76474
rect 6032 76424 6040 76474
rect 5714 76406 6040 76424
rect 5714 76332 6040 76350
rect 5714 76282 6015 76332
rect 6032 76282 6040 76332
rect 5714 76264 6040 76282
rect 5714 76190 6040 76208
rect 5714 76140 6015 76190
rect 6032 76140 6040 76190
rect 5714 76122 6040 76140
rect 5714 76048 6040 76066
rect 5714 75998 6015 76048
rect 6032 75998 6040 76048
rect 5714 75980 6040 75998
rect 5714 75906 6040 75924
rect 5714 75856 6015 75906
rect 6032 75856 6040 75906
rect 5714 75838 6040 75856
rect 5714 75764 6040 75782
rect 5714 75714 6015 75764
rect 6032 75714 6040 75764
rect 5714 75696 6040 75714
rect 5714 75622 6040 75640
rect 5714 75572 6015 75622
rect 6032 75572 6040 75622
rect 5714 75554 6040 75572
rect 5714 75480 6040 75498
rect 5714 75430 6015 75480
rect 6032 75430 6040 75480
rect 5714 75412 6040 75430
rect 5714 75338 6040 75356
rect 5714 75288 6015 75338
rect 6032 75288 6040 75338
rect 5714 75270 6040 75288
rect 5714 75196 6040 75214
rect 5714 75146 6015 75196
rect 6032 75146 6040 75196
rect 5714 75128 6040 75146
rect 5714 75054 6040 75072
rect 5714 75004 6015 75054
rect 6032 75004 6040 75054
rect 5714 74986 6040 75004
rect 5714 74912 6040 74930
rect 5714 74862 6015 74912
rect 6032 74862 6040 74912
rect 5714 74844 6040 74862
rect 5714 74770 6040 74788
rect 5714 74720 6015 74770
rect 6032 74720 6040 74770
rect 5714 74702 6040 74720
rect 5714 74628 6040 74646
rect 5714 74578 6015 74628
rect 6032 74578 6040 74628
rect 5714 74560 6040 74578
rect 5714 74486 6040 74504
rect 5714 74436 6015 74486
rect 6032 74436 6040 74486
rect 5714 74418 6040 74436
rect 5714 74344 6040 74362
rect 5714 74294 6015 74344
rect 6032 74294 6040 74344
rect 5714 74276 6040 74294
rect 5714 74202 6040 74220
rect 5714 74152 6015 74202
rect 6032 74152 6040 74202
rect 5714 74134 6040 74152
rect 5714 74060 6040 74078
rect 5714 74010 6015 74060
rect 6032 74010 6040 74060
rect 5714 73992 6040 74010
rect 5714 73918 6040 73936
rect 5714 73868 6015 73918
rect 6032 73868 6040 73918
rect 5714 73850 6040 73868
rect 5714 73776 6040 73794
rect 5714 73726 6015 73776
rect 6032 73726 6040 73776
rect 5714 73708 6040 73726
rect 5714 73634 6040 73652
rect 5714 73584 6015 73634
rect 6032 73584 6040 73634
rect 5714 73566 6040 73584
rect 5714 73492 6040 73510
rect 5714 73442 6015 73492
rect 6032 73442 6040 73492
rect 5714 73424 6040 73442
rect 5714 73350 6040 73368
rect 5714 73300 6015 73350
rect 6032 73300 6040 73350
rect 5714 73282 6040 73300
rect 5714 73208 6040 73226
rect 5714 73158 6015 73208
rect 6032 73158 6040 73208
rect 5714 73140 6040 73158
rect 5714 73066 6040 73084
rect 5714 73016 6015 73066
rect 6032 73016 6040 73066
rect 5714 72998 6040 73016
rect 5714 72924 6040 72942
rect 5714 72874 6015 72924
rect 6032 72874 6040 72924
rect 5714 72856 6040 72874
rect 5714 72782 6040 72800
rect 5714 72732 6015 72782
rect 6032 72732 6040 72782
rect 5714 72714 6040 72732
rect 5714 72640 6040 72658
rect 5714 72590 6015 72640
rect 6032 72590 6040 72640
rect 5714 72572 6040 72590
rect 5714 72498 6040 72516
rect 5714 72448 6015 72498
rect 6032 72448 6040 72498
rect 5714 72430 6040 72448
rect 5714 72356 6040 72374
rect 5714 72306 6015 72356
rect 6032 72306 6040 72356
rect 5714 72288 6040 72306
rect 5714 72214 6040 72232
rect 5714 72164 6015 72214
rect 6032 72164 6040 72214
rect 5714 72146 6040 72164
rect 5714 72072 6040 72090
rect 5714 72022 6015 72072
rect 6032 72022 6040 72072
rect 5714 72004 6040 72022
rect 5714 71930 6040 71948
rect 5714 71880 6015 71930
rect 6032 71880 6040 71930
rect 5714 71862 6040 71880
rect 5714 71788 6040 71806
rect 5714 71738 6015 71788
rect 6032 71738 6040 71788
rect 5714 71720 6040 71738
rect 5714 71646 6040 71664
rect 5714 71596 6015 71646
rect 6032 71596 6040 71646
rect 5714 71578 6040 71596
rect 5714 71504 6040 71522
rect 5714 71454 6015 71504
rect 6032 71454 6040 71504
rect 5714 71436 6040 71454
rect 5714 71362 6040 71380
rect 5714 71312 6015 71362
rect 6032 71312 6040 71362
rect 5714 71294 6040 71312
rect 5714 71220 6040 71238
rect 5714 71170 6015 71220
rect 6032 71170 6040 71220
rect 5714 71152 6040 71170
rect 5714 71078 6040 71096
rect 5714 71028 6015 71078
rect 6032 71028 6040 71078
rect 5714 71010 6040 71028
rect 5714 70936 6040 70954
rect 5714 70886 6015 70936
rect 6032 70886 6040 70936
rect 5714 70868 6040 70886
rect 5714 70794 6040 70812
rect 5714 70744 6015 70794
rect 6032 70744 6040 70794
rect 5714 70726 6040 70744
rect 5714 70652 6040 70670
rect 5714 70602 6015 70652
rect 6032 70602 6040 70652
rect 5714 70584 6040 70602
rect 5714 70510 6040 70528
rect 5714 70460 6015 70510
rect 6032 70460 6040 70510
rect 5714 70442 6040 70460
rect 5714 70368 6040 70386
rect 5714 70318 6015 70368
rect 6032 70318 6040 70368
rect 5714 70300 6040 70318
rect 5714 70226 6040 70244
rect 5714 70176 6015 70226
rect 6032 70176 6040 70226
rect 5714 70158 6040 70176
rect 5714 70084 6040 70102
rect 5714 70034 6015 70084
rect 6032 70034 6040 70084
rect 5714 70016 6040 70034
rect 5714 69942 6040 69960
rect 5714 69892 6015 69942
rect 6032 69892 6040 69942
rect 5714 69874 6040 69892
rect 5714 69800 6040 69818
rect 5714 69750 6015 69800
rect 6032 69750 6040 69800
rect 5714 69732 6040 69750
rect 5714 69658 6040 69676
rect 5714 69608 6015 69658
rect 6032 69608 6040 69658
rect 5714 69590 6040 69608
rect 5714 69516 6040 69534
rect 5714 69466 6015 69516
rect 6032 69466 6040 69516
rect 5714 69448 6040 69466
rect 5714 69374 6040 69392
rect 5714 69324 6015 69374
rect 6032 69324 6040 69374
rect 5714 69306 6040 69324
rect 5714 69232 6040 69250
rect 5714 69182 6015 69232
rect 6032 69182 6040 69232
rect 5714 69164 6040 69182
rect 5714 69090 6040 69108
rect 5714 69040 6015 69090
rect 6032 69040 6040 69090
rect 5714 69022 6040 69040
rect 5714 68948 6040 68966
rect 5714 68898 6015 68948
rect 6032 68898 6040 68948
rect 5714 68880 6040 68898
rect 5714 68806 6040 68824
rect 5714 68756 6015 68806
rect 6032 68756 6040 68806
rect 5714 68738 6040 68756
rect 5714 68664 6040 68682
rect 5714 68614 6015 68664
rect 6032 68614 6040 68664
rect 5714 68596 6040 68614
rect 5714 68522 6040 68540
rect 5714 68472 6015 68522
rect 6032 68472 6040 68522
rect 5714 68454 6040 68472
rect 5714 68380 6040 68398
rect 5714 68330 6015 68380
rect 6032 68330 6040 68380
rect 5714 68312 6040 68330
rect 5714 68238 6040 68256
rect 5714 68188 6015 68238
rect 6032 68188 6040 68238
rect 5714 68170 6040 68188
rect 5714 68096 6040 68114
rect 5714 68046 6015 68096
rect 6032 68046 6040 68096
rect 5714 68028 6040 68046
rect 5714 67954 6040 67972
rect 5714 67904 6015 67954
rect 6032 67904 6040 67954
rect 5714 67886 6040 67904
rect 5714 67812 6040 67830
rect 5714 67762 6015 67812
rect 6032 67762 6040 67812
rect 5714 67744 6040 67762
rect 5714 67670 6040 67688
rect 5714 67620 6015 67670
rect 6032 67620 6040 67670
rect 5714 67602 6040 67620
rect 5714 67528 6040 67546
rect 5714 67478 6015 67528
rect 6032 67478 6040 67528
rect 5714 67460 6040 67478
rect 5714 67386 6040 67404
rect 5714 67336 6015 67386
rect 6032 67336 6040 67386
rect 5714 67318 6040 67336
rect 5714 67244 6040 67262
rect 5714 67194 6015 67244
rect 6032 67194 6040 67244
rect 5714 67176 6040 67194
rect 5714 67102 6040 67120
rect 5714 67052 6015 67102
rect 6032 67052 6040 67102
rect 5714 67034 6040 67052
rect 5714 66960 6040 66978
rect 5714 66910 6015 66960
rect 6032 66910 6040 66960
rect 5714 66892 6040 66910
rect 5714 66818 6040 66836
rect 5714 66768 6015 66818
rect 6032 66768 6040 66818
rect 5714 66750 6040 66768
rect 5714 66676 6040 66694
rect 5714 66626 6015 66676
rect 6032 66626 6040 66676
rect 5714 66608 6040 66626
rect 5714 66534 6040 66552
rect 5714 66484 6015 66534
rect 6032 66484 6040 66534
rect 5714 66466 6040 66484
rect 5714 66392 6040 66410
rect 5714 66342 6015 66392
rect 6032 66342 6040 66392
rect 5714 66324 6040 66342
rect 5714 66250 6040 66268
rect 5714 66200 6015 66250
rect 6032 66200 6040 66250
rect 5714 66182 6040 66200
rect 5714 66108 6040 66126
rect 5714 66058 6015 66108
rect 6032 66058 6040 66108
rect 5714 66040 6040 66058
rect 5714 65966 6040 65984
rect 5714 65916 6015 65966
rect 6032 65916 6040 65966
rect 5714 65898 6040 65916
rect 5714 65824 6040 65842
rect 5714 65774 6015 65824
rect 6032 65774 6040 65824
rect 5714 65756 6040 65774
rect 5714 65682 6040 65700
rect 5714 65632 6015 65682
rect 6032 65632 6040 65682
rect 5714 65614 6040 65632
rect 5714 65540 6040 65558
rect 5714 65490 6015 65540
rect 6032 65490 6040 65540
rect 5714 65472 6040 65490
rect 5714 65398 6040 65416
rect 5714 65348 6015 65398
rect 6032 65348 6040 65398
rect 5714 65330 6040 65348
rect 5714 65256 6040 65274
rect 5714 65206 6015 65256
rect 6032 65206 6040 65256
rect 5714 65188 6040 65206
rect 5714 65114 6040 65132
rect 5714 65064 6015 65114
rect 6032 65064 6040 65114
rect 5714 65046 6040 65064
rect 5714 64972 6040 64990
rect 5714 64922 6015 64972
rect 6032 64922 6040 64972
rect 5714 64904 6040 64922
rect 5714 64830 6040 64848
rect 5714 64780 6015 64830
rect 6032 64780 6040 64830
rect 5714 64762 6040 64780
rect 5714 64688 6040 64706
rect 5714 64638 6015 64688
rect 6032 64638 6040 64688
rect 5714 64620 6040 64638
rect 5714 64546 6040 64564
rect 5714 64496 6015 64546
rect 6032 64496 6040 64546
rect 5714 64478 6040 64496
rect 5714 64404 6040 64422
rect 5714 64354 6015 64404
rect 6032 64354 6040 64404
rect 5714 64336 6040 64354
rect 5714 64262 6040 64280
rect 5714 64212 6015 64262
rect 6032 64212 6040 64262
rect 5714 64194 6040 64212
rect 5714 64120 6040 64138
rect 5714 64070 6015 64120
rect 6032 64070 6040 64120
rect 5714 64052 6040 64070
rect 5714 63978 6040 63996
rect 5714 63928 6015 63978
rect 6032 63928 6040 63978
rect 5714 63910 6040 63928
rect 5714 63836 6040 63854
rect 5714 63786 6015 63836
rect 6032 63786 6040 63836
rect 5714 63768 6040 63786
rect 5714 63694 6040 63712
rect 5714 63644 6015 63694
rect 6032 63644 6040 63694
rect 5714 63626 6040 63644
rect 5714 63552 6040 63570
rect 5714 63502 6015 63552
rect 6032 63502 6040 63552
rect 5714 63484 6040 63502
rect 5714 63410 6040 63428
rect 5714 63360 6015 63410
rect 6032 63360 6040 63410
rect 5714 63342 6040 63360
rect 5714 63268 6040 63286
rect 5714 63218 6015 63268
rect 6032 63218 6040 63268
rect 5714 63200 6040 63218
rect 5714 63126 6040 63144
rect 5714 63076 6015 63126
rect 6032 63076 6040 63126
rect 5714 63058 6040 63076
rect 5714 62984 6040 63002
rect 5714 62934 6015 62984
rect 6032 62934 6040 62984
rect 5714 62916 6040 62934
rect 5714 62842 6040 62860
rect 5714 62792 6015 62842
rect 6032 62792 6040 62842
rect 5714 62774 6040 62792
rect 5714 62700 6040 62718
rect 5714 62650 6015 62700
rect 6032 62650 6040 62700
rect 5714 62632 6040 62650
rect 5714 62558 6040 62576
rect 5714 62508 6015 62558
rect 6032 62508 6040 62558
rect 5714 62490 6040 62508
rect 5714 62416 6040 62434
rect 5714 62366 6015 62416
rect 6032 62366 6040 62416
rect 5714 62348 6040 62366
rect 5714 62274 6040 62292
rect 5714 62224 6015 62274
rect 6032 62224 6040 62274
rect 5714 62206 6040 62224
rect 5714 62132 6040 62150
rect 5714 62082 6015 62132
rect 6032 62082 6040 62132
rect 5714 62064 6040 62082
rect 5714 61990 6040 62008
rect 5714 61940 6015 61990
rect 6032 61940 6040 61990
rect 5714 61922 6040 61940
rect 5714 61848 6040 61866
rect 5714 61798 6015 61848
rect 6032 61798 6040 61848
rect 5714 61780 6040 61798
rect 5714 61706 6040 61724
rect 5714 61656 6015 61706
rect 6032 61656 6040 61706
rect 5714 61638 6040 61656
rect 5714 61564 6040 61582
rect 5714 61514 6015 61564
rect 6032 61514 6040 61564
rect 5714 61496 6040 61514
rect 5714 61422 6040 61440
rect 5714 61372 6015 61422
rect 6032 61372 6040 61422
rect 5714 61354 6040 61372
rect 5714 61280 6040 61298
rect 5714 61230 6015 61280
rect 6032 61230 6040 61280
rect 5714 61212 6040 61230
rect 5714 61138 6040 61156
rect 5714 61088 6015 61138
rect 6032 61088 6040 61138
rect 5714 61070 6040 61088
rect 5714 60996 6040 61014
rect 5714 60946 6015 60996
rect 6032 60946 6040 60996
rect 5714 60928 6040 60946
rect 5714 60854 6040 60872
rect 5714 60804 6015 60854
rect 6032 60804 6040 60854
rect 5714 60786 6040 60804
rect 5714 60712 6040 60730
rect 5714 60662 6015 60712
rect 6032 60662 6040 60712
rect 5714 60644 6040 60662
rect 5714 60570 6040 60588
rect 5714 60520 6015 60570
rect 6032 60520 6040 60570
rect 5714 60502 6040 60520
rect 5714 60428 6040 60446
rect 5714 60378 6015 60428
rect 6032 60378 6040 60428
rect 5714 60360 6040 60378
rect 5714 60286 6040 60304
rect 5714 60236 6015 60286
rect 6032 60236 6040 60286
rect 5714 60218 6040 60236
rect 5714 60144 6040 60162
rect 5714 60094 6015 60144
rect 6032 60094 6040 60144
rect 5714 60076 6040 60094
rect 5714 60002 6040 60020
rect 5714 59952 6015 60002
rect 6032 59952 6040 60002
rect 5714 59934 6040 59952
rect 5714 59860 6040 59878
rect 5714 59810 6015 59860
rect 6032 59810 6040 59860
rect 5714 59792 6040 59810
rect 5714 59718 6040 59736
rect 5714 59668 6015 59718
rect 6032 59668 6040 59718
rect 5714 59650 6040 59668
rect 5714 59576 6040 59594
rect 5714 59526 6015 59576
rect 6032 59526 6040 59576
rect 5714 59508 6040 59526
rect 5714 59434 6040 59452
rect 5714 59384 6015 59434
rect 6032 59384 6040 59434
rect 5714 59366 6040 59384
rect 5714 59292 6040 59310
rect 5714 59242 6015 59292
rect 6032 59242 6040 59292
rect 5714 59224 6040 59242
rect 5714 59150 6040 59168
rect 5714 59100 6015 59150
rect 6032 59100 6040 59150
rect 5714 59082 6040 59100
rect 5714 59008 6040 59026
rect 5714 58958 6015 59008
rect 6032 58958 6040 59008
rect 5714 58940 6040 58958
rect 5714 58866 6040 58884
rect 5714 58816 6015 58866
rect 6032 58816 6040 58866
rect 5714 58798 6040 58816
rect 5714 58724 6040 58742
rect 5714 58674 6015 58724
rect 6032 58674 6040 58724
rect 5714 58656 6040 58674
rect 5714 58582 6040 58600
rect 5714 58532 6015 58582
rect 6032 58532 6040 58582
rect 5714 58514 6040 58532
rect 5714 58440 6040 58458
rect 5714 58390 6015 58440
rect 6032 58390 6040 58440
rect 5714 58372 6040 58390
rect 5714 58298 6040 58316
rect 5714 58248 6015 58298
rect 6032 58248 6040 58298
rect 5714 58230 6040 58248
rect 5714 58156 6040 58174
rect 5714 58106 6015 58156
rect 6032 58106 6040 58156
rect 5714 58088 6040 58106
rect 5714 58014 6040 58032
rect 5714 57964 6015 58014
rect 6032 57964 6040 58014
rect 5714 57946 6040 57964
rect 5714 57872 6040 57890
rect 5714 57822 6015 57872
rect 6032 57822 6040 57872
rect 5714 57804 6040 57822
rect 5714 57730 6040 57748
rect 5714 57680 6015 57730
rect 6032 57680 6040 57730
rect 5714 57662 6040 57680
rect 5714 57588 6040 57606
rect 5714 57538 6015 57588
rect 6032 57538 6040 57588
rect 5714 57520 6040 57538
rect 5714 57446 6040 57464
rect 5714 57396 6015 57446
rect 6032 57396 6040 57446
rect 5714 57378 6040 57396
rect 5714 57304 6040 57322
rect 5714 57254 6015 57304
rect 6032 57254 6040 57304
rect 5714 57236 6040 57254
rect 5714 57162 6040 57180
rect 5714 57112 6015 57162
rect 6032 57112 6040 57162
rect 5714 57094 6040 57112
rect 5714 57020 6040 57038
rect 5714 56970 6015 57020
rect 6032 56970 6040 57020
rect 5714 56952 6040 56970
rect 5714 56878 6040 56896
rect 5714 56828 6015 56878
rect 6032 56828 6040 56878
rect 5714 56810 6040 56828
rect 5714 56736 6040 56754
rect 5714 56686 6015 56736
rect 6032 56686 6040 56736
rect 5714 56668 6040 56686
rect 5714 56594 6040 56612
rect 5714 56544 6015 56594
rect 6032 56544 6040 56594
rect 5714 56526 6040 56544
rect 5714 56452 6040 56470
rect 5714 56402 6015 56452
rect 6032 56402 6040 56452
rect 5714 56384 6040 56402
rect 5714 56310 6040 56328
rect 5714 56260 6015 56310
rect 6032 56260 6040 56310
rect 5714 56242 6040 56260
rect 5714 56168 6040 56186
rect 5714 56118 6015 56168
rect 6032 56118 6040 56168
rect 5714 56100 6040 56118
rect 5714 56026 6040 56044
rect 5714 55976 6015 56026
rect 6032 55976 6040 56026
rect 5714 55958 6040 55976
rect 5714 55884 6040 55902
rect 5714 55834 6015 55884
rect 6032 55834 6040 55884
rect 5714 55816 6040 55834
rect 5714 55742 6040 55760
rect 5714 55692 6015 55742
rect 6032 55692 6040 55742
rect 5714 55674 6040 55692
rect 5714 55600 6040 55618
rect 5714 55550 6015 55600
rect 6032 55550 6040 55600
rect 5714 55532 6040 55550
rect 5714 55458 6040 55476
rect 5714 55408 6015 55458
rect 6032 55408 6040 55458
rect 5714 55390 6040 55408
rect 5714 55316 6040 55334
rect 5714 55266 6015 55316
rect 6032 55266 6040 55316
rect 5714 55248 6040 55266
rect 5714 55174 6040 55192
rect 5714 55124 6015 55174
rect 6032 55124 6040 55174
rect 5714 55106 6040 55124
rect 5714 55032 6040 55050
rect 5714 54982 6015 55032
rect 6032 54982 6040 55032
rect 5714 54964 6040 54982
rect 5714 54890 6040 54908
rect 5714 54840 6015 54890
rect 6032 54840 6040 54890
rect 5714 54822 6040 54840
rect 5714 54748 6040 54766
rect 5714 54698 6015 54748
rect 6032 54698 6040 54748
rect 5714 54680 6040 54698
rect 5714 54606 6040 54624
rect 5714 54556 6015 54606
rect 6032 54556 6040 54606
rect 5714 54538 6040 54556
rect 5714 54464 6040 54482
rect 5714 54414 6015 54464
rect 6032 54414 6040 54464
rect 5714 54396 6040 54414
rect 5714 54322 6040 54340
rect 5714 54272 6015 54322
rect 6032 54272 6040 54322
rect 5714 54254 6040 54272
rect 5714 54180 6040 54198
rect 5714 54130 6015 54180
rect 6032 54130 6040 54180
rect 5714 54112 6040 54130
rect 5714 54038 6040 54056
rect 5714 53988 6015 54038
rect 6032 53988 6040 54038
rect 5714 53970 6040 53988
rect 5714 53896 6040 53914
rect 5714 53846 6015 53896
rect 6032 53846 6040 53896
rect 5714 53828 6040 53846
rect 5714 53754 6040 53772
rect 5714 53704 6015 53754
rect 6032 53704 6040 53754
rect 5714 53686 6040 53704
rect 5714 53612 6040 53630
rect 5714 53562 6015 53612
rect 6032 53562 6040 53612
rect 5714 53544 6040 53562
rect 5714 53470 6040 53488
rect 5714 53420 6015 53470
rect 6032 53420 6040 53470
rect 5714 53402 6040 53420
rect 5714 53328 6040 53346
rect 5714 53278 6015 53328
rect 6032 53278 6040 53328
rect 5714 53260 6040 53278
rect 5714 53186 6040 53204
rect 5714 53136 6015 53186
rect 6032 53136 6040 53186
rect 5714 53118 6040 53136
rect 5714 53044 6040 53062
rect 5714 52994 6015 53044
rect 6032 52994 6040 53044
rect 5714 52976 6040 52994
rect 5714 52902 6040 52920
rect 5714 52852 6015 52902
rect 6032 52852 6040 52902
rect 5714 52834 6040 52852
rect 5714 52760 6040 52778
rect 5714 52710 6015 52760
rect 6032 52710 6040 52760
rect 5714 52692 6040 52710
rect 5714 52618 6040 52636
rect 5714 52568 6015 52618
rect 6032 52568 6040 52618
rect 5714 52550 6040 52568
rect 5714 52476 6040 52494
rect 5714 52426 6015 52476
rect 6032 52426 6040 52476
rect 5714 52408 6040 52426
rect 5714 52334 6040 52352
rect 5714 52284 6015 52334
rect 6032 52284 6040 52334
rect 5714 52266 6040 52284
rect 5714 52192 6040 52210
rect 5714 52142 6015 52192
rect 6032 52142 6040 52192
rect 5714 52124 6040 52142
rect 5714 52050 6040 52068
rect 5714 52000 6015 52050
rect 6032 52000 6040 52050
rect 5714 51982 6040 52000
rect 5714 51908 6040 51926
rect 5714 51858 6015 51908
rect 6032 51858 6040 51908
rect 5714 51840 6040 51858
rect 5714 51766 6040 51784
rect 5714 51716 6015 51766
rect 6032 51716 6040 51766
rect 5714 51698 6040 51716
rect 5714 51624 6040 51642
rect 5714 51574 6015 51624
rect 6032 51574 6040 51624
rect 5714 51556 6040 51574
rect 5714 51482 6040 51500
rect 5714 51432 6015 51482
rect 6032 51432 6040 51482
rect 5714 51414 6040 51432
rect 5714 51340 6040 51358
rect 5714 51290 6015 51340
rect 6032 51290 6040 51340
rect 5714 51272 6040 51290
rect 5714 51198 6040 51216
rect 5714 51148 6015 51198
rect 6032 51148 6040 51198
rect 5714 51130 6040 51148
rect 5714 51056 6040 51074
rect 5714 51006 6015 51056
rect 6032 51006 6040 51056
rect 5714 50988 6040 51006
rect 5714 50914 6040 50932
rect 5714 50864 6015 50914
rect 6032 50864 6040 50914
rect 5714 50846 6040 50864
rect 5714 50772 6040 50790
rect 5714 50722 6015 50772
rect 6032 50722 6040 50772
rect 5714 50704 6040 50722
rect 5714 50630 6040 50648
rect 5714 50580 6015 50630
rect 6032 50580 6040 50630
rect 5714 50562 6040 50580
rect 5714 50488 6040 50506
rect 5714 50438 6015 50488
rect 6032 50438 6040 50488
rect 5714 50420 6040 50438
rect 5714 50346 6040 50364
rect 5714 50296 6015 50346
rect 6032 50296 6040 50346
rect 5714 50278 6040 50296
rect 5714 50204 6040 50222
rect 5714 50154 6015 50204
rect 6032 50154 6040 50204
rect 5714 50136 6040 50154
rect 5714 50062 6040 50080
rect 5714 50012 6015 50062
rect 6032 50012 6040 50062
rect 5714 49994 6040 50012
rect 5714 49920 6040 49938
rect 5714 49870 6015 49920
rect 6032 49870 6040 49920
rect 5714 49852 6040 49870
rect 5714 49778 6040 49796
rect 5714 49728 6015 49778
rect 6032 49728 6040 49778
rect 5714 49710 6040 49728
rect 5714 49636 6040 49654
rect 5714 49586 6015 49636
rect 6032 49586 6040 49636
rect 5714 49568 6040 49586
rect 5714 49494 6040 49512
rect 5714 49444 6015 49494
rect 6032 49444 6040 49494
rect 5714 49426 6040 49444
rect 5714 49352 6040 49370
rect 5714 49302 6015 49352
rect 6032 49302 6040 49352
rect 5714 49284 6040 49302
rect 5714 49210 6040 49228
rect 5714 49160 6015 49210
rect 6032 49160 6040 49210
rect 5714 49142 6040 49160
rect 5714 49068 6040 49086
rect 5714 49018 6015 49068
rect 6032 49018 6040 49068
rect 5714 49000 6040 49018
rect 5714 48926 6040 48944
rect 5714 48876 6015 48926
rect 6032 48876 6040 48926
rect 5714 48858 6040 48876
rect 5714 48784 6040 48802
rect 5714 48734 6015 48784
rect 6032 48734 6040 48784
rect 5714 48716 6040 48734
rect 5714 48642 6040 48660
rect 5714 48592 6015 48642
rect 6032 48592 6040 48642
rect 5714 48574 6040 48592
rect 5714 48500 6040 48518
rect 5714 48450 6015 48500
rect 6032 48450 6040 48500
rect 5714 48432 6040 48450
rect 5714 48358 6040 48376
rect 5714 48308 6015 48358
rect 6032 48308 6040 48358
rect 5714 48290 6040 48308
rect 5714 48216 6040 48234
rect 5714 48166 6015 48216
rect 6032 48166 6040 48216
rect 5714 48148 6040 48166
rect 5714 48074 6040 48092
rect 5714 48024 6015 48074
rect 6032 48024 6040 48074
rect 5714 48006 6040 48024
rect 5714 47932 6040 47950
rect 5714 47882 6015 47932
rect 6032 47882 6040 47932
rect 5714 47864 6040 47882
rect 5714 47790 6040 47808
rect 5714 47740 6015 47790
rect 6032 47740 6040 47790
rect 5714 47722 6040 47740
rect 5714 47648 6040 47666
rect 5714 47598 6015 47648
rect 6032 47598 6040 47648
rect 5714 47580 6040 47598
rect 5714 47506 6040 47524
rect 5714 47456 6015 47506
rect 6032 47456 6040 47506
rect 5714 47438 6040 47456
rect 5714 47364 6040 47382
rect 5714 47314 6015 47364
rect 6032 47314 6040 47364
rect 5714 47296 6040 47314
rect 5714 47222 6040 47240
rect 5714 47172 6015 47222
rect 6032 47172 6040 47222
rect 5714 47154 6040 47172
rect 5714 47080 6040 47098
rect 5714 47030 6015 47080
rect 6032 47030 6040 47080
rect 5714 47012 6040 47030
rect 5714 46938 6040 46956
rect 5714 46888 6015 46938
rect 6032 46888 6040 46938
rect 5714 46870 6040 46888
rect 5714 46796 6040 46814
rect 5714 46746 6015 46796
rect 6032 46746 6040 46796
rect 5714 46728 6040 46746
rect 5714 46654 6040 46672
rect 5714 46604 6015 46654
rect 6032 46604 6040 46654
rect 5714 46586 6040 46604
rect 5714 46512 6040 46530
rect 5714 46462 6015 46512
rect 6032 46462 6040 46512
rect 5714 46444 6040 46462
rect 5714 46370 6040 46388
rect 5714 46320 6015 46370
rect 6032 46320 6040 46370
rect 5714 46302 6040 46320
rect 5714 46228 6040 46246
rect 5714 46178 6015 46228
rect 6032 46178 6040 46228
rect 5714 46160 6040 46178
rect 5714 46086 6040 46104
rect 5714 46036 6015 46086
rect 6032 46036 6040 46086
rect 5714 46018 6040 46036
rect 5714 45944 6040 45962
rect 5714 45894 6015 45944
rect 6032 45894 6040 45944
rect 5714 45876 6040 45894
rect 5714 45802 6040 45820
rect 5714 45752 6015 45802
rect 6032 45752 6040 45802
rect 5714 45734 6040 45752
rect 5714 45660 6040 45678
rect 5714 45610 6015 45660
rect 6032 45610 6040 45660
rect 5714 45592 6040 45610
rect 5714 45518 6040 45536
rect 5714 45468 6015 45518
rect 6032 45468 6040 45518
rect 5714 45450 6040 45468
rect 5714 45376 6040 45394
rect 5714 45326 6015 45376
rect 6032 45326 6040 45376
rect 5714 45308 6040 45326
rect 5714 45234 6040 45252
rect 5714 45184 6015 45234
rect 6032 45184 6040 45234
rect 5714 45166 6040 45184
rect 5714 45092 6040 45110
rect 5714 45042 6015 45092
rect 6032 45042 6040 45092
rect 5714 45024 6040 45042
rect 5714 44950 6040 44968
rect 5714 44900 6015 44950
rect 6032 44900 6040 44950
rect 5714 44882 6040 44900
rect 5714 44808 6040 44826
rect 5714 44758 6015 44808
rect 6032 44758 6040 44808
rect 5714 44740 6040 44758
rect 5714 44666 6040 44684
rect 5714 44616 6015 44666
rect 6032 44616 6040 44666
rect 5714 44598 6040 44616
rect 5714 44524 6040 44542
rect 5714 44474 6015 44524
rect 6032 44474 6040 44524
rect 5714 44456 6040 44474
rect 5714 44382 6040 44400
rect 5714 44332 6015 44382
rect 6032 44332 6040 44382
rect 5714 44314 6040 44332
rect 5714 44240 6040 44258
rect 5714 44190 6015 44240
rect 6032 44190 6040 44240
rect 5714 44172 6040 44190
rect 5714 44098 6040 44116
rect 5714 44048 6015 44098
rect 6032 44048 6040 44098
rect 5714 44030 6040 44048
rect 5714 43956 6040 43974
rect 5714 43906 6015 43956
rect 6032 43906 6040 43956
rect 5714 43888 6040 43906
rect 5714 43814 6040 43832
rect 5714 43764 6015 43814
rect 6032 43764 6040 43814
rect 5714 43746 6040 43764
rect 5714 43672 6040 43690
rect 5714 43622 6015 43672
rect 6032 43622 6040 43672
rect 5714 43604 6040 43622
rect 5714 43530 6040 43548
rect 5714 43480 6015 43530
rect 6032 43480 6040 43530
rect 5714 43462 6040 43480
rect 5714 43388 6040 43406
rect 5714 43338 6015 43388
rect 6032 43338 6040 43388
rect 5714 43320 6040 43338
rect 5714 43246 6040 43264
rect 5714 43196 6015 43246
rect 6032 43196 6040 43246
rect 5714 43178 6040 43196
rect 5714 43104 6040 43122
rect 5714 43054 6015 43104
rect 6032 43054 6040 43104
rect 5714 43036 6040 43054
rect 5714 42962 6040 42980
rect 5714 42912 6015 42962
rect 6032 42912 6040 42962
rect 5714 42894 6040 42912
rect 5714 42820 6040 42838
rect 5714 42770 6015 42820
rect 6032 42770 6040 42820
rect 5714 42752 6040 42770
rect 5714 42678 6040 42696
rect 5714 42628 6015 42678
rect 6032 42628 6040 42678
rect 5714 42610 6040 42628
rect 5714 42536 6040 42554
rect 5714 42486 6015 42536
rect 6032 42486 6040 42536
rect 5714 42468 6040 42486
rect 5714 42394 6040 42412
rect 5714 42344 6015 42394
rect 6032 42344 6040 42394
rect 5714 42326 6040 42344
rect 5714 42252 6040 42270
rect 5714 42202 6015 42252
rect 6032 42202 6040 42252
rect 5714 42184 6040 42202
rect 5714 42110 6040 42128
rect 5714 42060 6015 42110
rect 6032 42060 6040 42110
rect 5714 42042 6040 42060
rect 5714 41968 6040 41986
rect 5714 41918 6015 41968
rect 6032 41918 6040 41968
rect 5714 41900 6040 41918
rect 5714 41826 6040 41844
rect 5714 41776 6015 41826
rect 6032 41776 6040 41826
rect 5714 41758 6040 41776
rect 5714 41684 6040 41702
rect 5714 41634 6015 41684
rect 6032 41634 6040 41684
rect 5714 41616 6040 41634
rect 5714 41542 6040 41560
rect 5714 41492 6015 41542
rect 6032 41492 6040 41542
rect 5714 41474 6040 41492
rect 5714 41400 6040 41418
rect 5714 41350 6015 41400
rect 6032 41350 6040 41400
rect 5714 41332 6040 41350
rect 5714 41258 6040 41276
rect 5714 41208 6015 41258
rect 6032 41208 6040 41258
rect 5714 41190 6040 41208
rect 5714 41116 6040 41134
rect 5714 41066 6015 41116
rect 6032 41066 6040 41116
rect 5714 41048 6040 41066
rect 5714 40974 6040 40992
rect 5714 40924 6015 40974
rect 6032 40924 6040 40974
rect 5714 40906 6040 40924
rect 5714 40832 6040 40850
rect 5714 40782 6015 40832
rect 6032 40782 6040 40832
rect 5714 40764 6040 40782
rect 5714 40690 6040 40708
rect 5714 40640 6015 40690
rect 6032 40640 6040 40690
rect 5714 40622 6040 40640
rect 5714 40548 6040 40566
rect 5714 40498 6015 40548
rect 6032 40498 6040 40548
rect 5714 40480 6040 40498
rect 5714 40406 6040 40424
rect 5714 40356 6015 40406
rect 6032 40356 6040 40406
rect 5714 40338 6040 40356
rect 5714 40264 6040 40282
rect 5714 40214 6015 40264
rect 6032 40214 6040 40264
rect 5714 40196 6040 40214
rect 5714 40122 6040 40140
rect 5714 40072 6015 40122
rect 6032 40072 6040 40122
rect 5714 40054 6040 40072
rect 5714 39980 6040 39998
rect 5714 39930 6015 39980
rect 6032 39930 6040 39980
rect 5714 39912 6040 39930
rect 5714 39838 6040 39856
rect 5714 39788 6015 39838
rect 6032 39788 6040 39838
rect 5714 39770 6040 39788
rect 5714 39696 6040 39714
rect 5714 39646 6015 39696
rect 6032 39646 6040 39696
rect 5714 39628 6040 39646
rect 5714 39554 6040 39572
rect 5714 39504 6015 39554
rect 6032 39504 6040 39554
rect 5714 39486 6040 39504
rect 5714 39412 6040 39430
rect 5714 39362 6015 39412
rect 6032 39362 6040 39412
rect 5714 39344 6040 39362
rect 5714 39270 6040 39288
rect 5714 39220 6015 39270
rect 6032 39220 6040 39270
rect 5714 39202 6040 39220
rect 5714 39128 6040 39146
rect 5714 39078 6015 39128
rect 6032 39078 6040 39128
rect 5714 39060 6040 39078
rect 5714 38986 6040 39004
rect 5714 38936 6015 38986
rect 6032 38936 6040 38986
rect 5714 38918 6040 38936
rect 5714 38844 6040 38862
rect 5714 38794 6015 38844
rect 6032 38794 6040 38844
rect 5714 38776 6040 38794
rect 5714 38702 6040 38720
rect 5714 38652 6015 38702
rect 6032 38652 6040 38702
rect 5714 38634 6040 38652
rect 5714 38560 6040 38578
rect 5714 38510 6015 38560
rect 6032 38510 6040 38560
rect 5714 38492 6040 38510
rect 5714 38418 6040 38436
rect 5714 38368 6015 38418
rect 6032 38368 6040 38418
rect 5714 38350 6040 38368
rect 5714 38276 6040 38294
rect 5714 38226 6015 38276
rect 6032 38226 6040 38276
rect 5714 38208 6040 38226
rect 5714 38134 6040 38152
rect 5714 38084 6015 38134
rect 6032 38084 6040 38134
rect 5714 38066 6040 38084
rect 5714 37992 6040 38010
rect 5714 37942 6015 37992
rect 6032 37942 6040 37992
rect 5714 37924 6040 37942
rect 5714 37850 6040 37868
rect 5714 37800 6015 37850
rect 6032 37800 6040 37850
rect 5714 37782 6040 37800
rect 5714 37708 6040 37726
rect 5714 37658 6015 37708
rect 6032 37658 6040 37708
rect 5714 37640 6040 37658
rect 5714 37566 6040 37584
rect 5714 37516 6015 37566
rect 6032 37516 6040 37566
rect 5714 37498 6040 37516
rect 5714 37424 6040 37442
rect 5714 37374 6015 37424
rect 6032 37374 6040 37424
rect 5714 37356 6040 37374
rect 5714 37282 6040 37300
rect 5714 37232 6015 37282
rect 6032 37232 6040 37282
rect 5714 37214 6040 37232
rect 5714 37140 6040 37158
rect 5714 37090 6015 37140
rect 6032 37090 6040 37140
rect 5714 37072 6040 37090
rect 5714 36998 6040 37016
rect 5714 36948 6015 36998
rect 6032 36948 6040 36998
rect 5714 36930 6040 36948
rect 5714 36856 6040 36874
rect 5714 36806 6015 36856
rect 6032 36806 6040 36856
rect 5714 36788 6040 36806
rect 5714 36714 6040 36732
rect 5714 36664 6015 36714
rect 6032 36664 6040 36714
rect 5714 36646 6040 36664
rect 5714 36572 6040 36590
rect 5714 36522 6015 36572
rect 6032 36522 6040 36572
rect 5714 36504 6040 36522
rect 5714 36430 6040 36448
rect 5714 36380 6015 36430
rect 6032 36380 6040 36430
rect 5714 36362 6040 36380
rect 5714 36288 6040 36306
rect 5714 36238 6015 36288
rect 6032 36238 6040 36288
rect 5714 36220 6040 36238
rect 5714 36146 6040 36164
rect 5714 36096 6015 36146
rect 6032 36096 6040 36146
rect 5714 36078 6040 36096
rect 5714 36004 6040 36022
rect 5714 35954 6015 36004
rect 6032 35954 6040 36004
rect 5714 35936 6040 35954
rect 5714 35862 6040 35880
rect 5714 35812 6015 35862
rect 6032 35812 6040 35862
rect 5714 35794 6040 35812
rect 5714 35720 6040 35738
rect 5714 35670 6015 35720
rect 6032 35670 6040 35720
rect 5714 35652 6040 35670
rect 5714 35578 6040 35596
rect 5714 35528 6015 35578
rect 6032 35528 6040 35578
rect 5714 35510 6040 35528
rect 5714 35436 6040 35454
rect 5714 35386 6015 35436
rect 6032 35386 6040 35436
rect 5714 35368 6040 35386
rect 5714 35294 6040 35312
rect 5714 35244 6015 35294
rect 6032 35244 6040 35294
rect 5714 35226 6040 35244
rect 5714 35152 6040 35170
rect 5714 35102 6015 35152
rect 6032 35102 6040 35152
rect 5714 35084 6040 35102
rect 5714 35010 6040 35028
rect 5714 34960 6015 35010
rect 6032 34960 6040 35010
rect 5714 34942 6040 34960
rect 5714 34868 6040 34886
rect 5714 34818 6015 34868
rect 6032 34818 6040 34868
rect 5714 34800 6040 34818
rect 5714 34726 6040 34744
rect 5714 34676 6015 34726
rect 6032 34676 6040 34726
rect 5714 34658 6040 34676
rect 5714 34584 6040 34602
rect 5714 34534 6015 34584
rect 6032 34534 6040 34584
rect 5714 34516 6040 34534
rect 5714 34442 6040 34460
rect 5714 34392 6015 34442
rect 6032 34392 6040 34442
rect 5714 34374 6040 34392
rect 5714 34300 6040 34318
rect 5714 34250 6015 34300
rect 6032 34250 6040 34300
rect 5714 34232 6040 34250
rect 5714 34158 6040 34176
rect 5714 34108 6015 34158
rect 6032 34108 6040 34158
rect 5714 34090 6040 34108
rect 5714 34016 6040 34034
rect 5714 33966 6015 34016
rect 6032 33966 6040 34016
rect 5714 33948 6040 33966
rect 5714 33874 6040 33892
rect 5714 33824 6015 33874
rect 6032 33824 6040 33874
rect 5714 33806 6040 33824
rect 5714 33732 6040 33750
rect 5714 33682 6015 33732
rect 6032 33682 6040 33732
rect 5714 33664 6040 33682
rect 5714 33590 6040 33608
rect 5714 33540 6015 33590
rect 6032 33540 6040 33590
rect 5714 33522 6040 33540
rect 5714 33448 6040 33466
rect 5714 33398 6015 33448
rect 6032 33398 6040 33448
rect 5714 33380 6040 33398
rect 5714 33306 6040 33324
rect 5714 33256 6015 33306
rect 6032 33256 6040 33306
rect 5714 33238 6040 33256
rect 5714 33164 6040 33182
rect 5714 33114 6015 33164
rect 6032 33114 6040 33164
rect 5714 33096 6040 33114
rect 5714 33022 6040 33040
rect 5714 32972 6015 33022
rect 6032 32972 6040 33022
rect 5714 32954 6040 32972
rect 5714 32880 6040 32898
rect 5714 32830 6015 32880
rect 6032 32830 6040 32880
rect 5714 32812 6040 32830
rect 5714 32738 6040 32756
rect 5714 32688 6015 32738
rect 6032 32688 6040 32738
rect 5714 32670 6040 32688
rect 5714 32596 6040 32614
rect 5714 32546 6015 32596
rect 6032 32546 6040 32596
rect 5714 32528 6040 32546
rect 5714 32454 6040 32472
rect 5714 32404 6015 32454
rect 6032 32404 6040 32454
rect 5714 32386 6040 32404
rect 5714 32312 6040 32330
rect 5714 32262 6015 32312
rect 6032 32262 6040 32312
rect 5714 32244 6040 32262
rect 5714 32170 6040 32188
rect 5714 32120 6015 32170
rect 6032 32120 6040 32170
rect 5714 32102 6040 32120
rect 5714 32028 6040 32046
rect 5714 31978 6015 32028
rect 6032 31978 6040 32028
rect 5714 31960 6040 31978
rect 5714 31886 6040 31904
rect 5714 31836 6015 31886
rect 6032 31836 6040 31886
rect 5714 31818 6040 31836
rect 5714 31744 6040 31762
rect 5714 31694 6015 31744
rect 6032 31694 6040 31744
rect 5714 31676 6040 31694
rect 5714 31602 6040 31620
rect 5714 31552 6015 31602
rect 6032 31552 6040 31602
rect 5714 31534 6040 31552
rect 5714 31460 6040 31478
rect 5714 31410 6015 31460
rect 6032 31410 6040 31460
rect 5714 31392 6040 31410
rect 5714 31318 6040 31336
rect 5714 31268 6015 31318
rect 6032 31268 6040 31318
rect 5714 31250 6040 31268
rect 5714 31176 6040 31194
rect 5714 31126 6015 31176
rect 6032 31126 6040 31176
rect 5714 31108 6040 31126
rect 5714 31034 6040 31052
rect 5714 30984 6015 31034
rect 6032 30984 6040 31034
rect 5714 30966 6040 30984
rect 5714 30892 6040 30910
rect 5714 30842 6015 30892
rect 6032 30842 6040 30892
rect 5714 30824 6040 30842
rect 5714 30750 6040 30768
rect 5714 30700 6015 30750
rect 6032 30700 6040 30750
rect 5714 30682 6040 30700
rect 5714 30608 6040 30626
rect 5714 30558 6015 30608
rect 6032 30558 6040 30608
rect 5714 30540 6040 30558
rect 5714 30466 6040 30484
rect 5714 30416 6015 30466
rect 6032 30416 6040 30466
rect 5714 30398 6040 30416
rect 5714 30324 6040 30342
rect 5714 30274 6015 30324
rect 6032 30274 6040 30324
rect 5714 30256 6040 30274
rect 5714 30182 6040 30200
rect 5714 30132 6015 30182
rect 6032 30132 6040 30182
rect 5714 30114 6040 30132
rect 5714 30040 6040 30058
rect 5714 29990 6015 30040
rect 6032 29990 6040 30040
rect 5714 29972 6040 29990
rect 5714 29898 6040 29916
rect 5714 29848 6015 29898
rect 6032 29848 6040 29898
rect 5714 29830 6040 29848
rect 5714 29756 6040 29774
rect 5714 29706 6015 29756
rect 6032 29706 6040 29756
rect 5714 29688 6040 29706
rect 5714 29614 6040 29632
rect 5714 29564 6015 29614
rect 6032 29564 6040 29614
rect 5714 29546 6040 29564
rect 5714 29472 6040 29490
rect 5714 29422 6015 29472
rect 6032 29422 6040 29472
rect 5714 29404 6040 29422
rect 5714 29330 6040 29348
rect 5714 29280 6015 29330
rect 6032 29280 6040 29330
rect 5714 29262 6040 29280
rect 5714 29188 6040 29206
rect 5714 29138 6015 29188
rect 6032 29138 6040 29188
rect 5714 29120 6040 29138
rect 5714 29046 6040 29064
rect 5714 28996 6015 29046
rect 6032 28996 6040 29046
rect 5714 28978 6040 28996
rect 5714 28904 6040 28922
rect 5714 28854 6015 28904
rect 6032 28854 6040 28904
rect 5714 28836 6040 28854
rect 5714 28762 6040 28780
rect 5714 28712 6015 28762
rect 6032 28712 6040 28762
rect 5714 28694 6040 28712
rect 5714 28620 6040 28638
rect 5714 28570 6015 28620
rect 6032 28570 6040 28620
rect 5714 28552 6040 28570
rect 5714 28478 6040 28496
rect 5714 28428 6015 28478
rect 6032 28428 6040 28478
rect 5714 28410 6040 28428
rect 5714 28336 6040 28354
rect 5714 28286 6015 28336
rect 6032 28286 6040 28336
rect 5714 28268 6040 28286
rect 5714 28194 6040 28212
rect 5714 28144 6015 28194
rect 6032 28144 6040 28194
rect 5714 28126 6040 28144
rect 5714 28052 6040 28070
rect 5714 28002 6015 28052
rect 6032 28002 6040 28052
rect 5714 27984 6040 28002
rect 5714 27910 6040 27928
rect 5714 27860 6015 27910
rect 6032 27860 6040 27910
rect 5714 27842 6040 27860
rect 5714 27768 6040 27786
rect 5714 27718 6015 27768
rect 6032 27718 6040 27768
rect 5714 27700 6040 27718
rect 5714 27626 6040 27644
rect 5714 27576 6015 27626
rect 6032 27576 6040 27626
rect 5714 27558 6040 27576
rect 5714 27484 6040 27502
rect 5714 27434 6015 27484
rect 6032 27434 6040 27484
rect 5714 27416 6040 27434
rect 5714 27342 6040 27360
rect 5714 27292 6015 27342
rect 6032 27292 6040 27342
rect 5714 27274 6040 27292
rect 5714 27200 6040 27218
rect 5714 27150 6015 27200
rect 6032 27150 6040 27200
rect 5714 27132 6040 27150
rect 5714 27058 6040 27076
rect 5714 27008 6015 27058
rect 6032 27008 6040 27058
rect 5714 26990 6040 27008
rect 5714 26916 6040 26934
rect 5714 26866 6015 26916
rect 6032 26866 6040 26916
rect 5714 26848 6040 26866
rect 5714 26774 6040 26792
rect 5714 26724 6015 26774
rect 6032 26724 6040 26774
rect 5714 26706 6040 26724
rect 5714 26632 6040 26650
rect 5714 26582 6015 26632
rect 6032 26582 6040 26632
rect 5714 26564 6040 26582
rect 5714 26490 6040 26508
rect 5714 26440 6015 26490
rect 6032 26440 6040 26490
rect 5714 26422 6040 26440
rect 5714 26348 6040 26366
rect 5714 26298 6015 26348
rect 6032 26298 6040 26348
rect 5714 26280 6040 26298
rect 5714 26206 6040 26224
rect 5714 26156 6015 26206
rect 6032 26156 6040 26206
rect 5714 26138 6040 26156
rect 5714 26064 6040 26082
rect 5714 26014 6015 26064
rect 6032 26014 6040 26064
rect 5714 25996 6040 26014
rect 5714 25922 6040 25940
rect 5714 25872 6015 25922
rect 6032 25872 6040 25922
rect 5714 25854 6040 25872
rect 5714 25780 6040 25798
rect 5714 25730 6015 25780
rect 6032 25730 6040 25780
rect 5714 25712 6040 25730
rect 5714 25638 6040 25656
rect 5714 25588 6015 25638
rect 6032 25588 6040 25638
rect 5714 25570 6040 25588
rect 5714 25496 6040 25514
rect 5714 25446 6015 25496
rect 6032 25446 6040 25496
rect 5714 25428 6040 25446
rect 5714 25354 6040 25372
rect 5714 25304 6015 25354
rect 6032 25304 6040 25354
rect 5714 25286 6040 25304
rect 5714 25212 6040 25230
rect 5714 25162 6015 25212
rect 6032 25162 6040 25212
rect 5714 25144 6040 25162
rect 5714 25070 6040 25088
rect 5714 25020 6015 25070
rect 6032 25020 6040 25070
rect 5714 25002 6040 25020
rect 5714 24928 6040 24946
rect 5714 24878 6015 24928
rect 6032 24878 6040 24928
rect 5714 24860 6040 24878
rect 5714 24786 6040 24804
rect 5714 24736 6015 24786
rect 6032 24736 6040 24786
rect 5714 24718 6040 24736
rect 5714 24644 6040 24662
rect 5714 24594 6015 24644
rect 6032 24594 6040 24644
rect 5714 24576 6040 24594
rect 5714 24502 6040 24520
rect 5714 24452 6015 24502
rect 6032 24452 6040 24502
rect 5714 24434 6040 24452
rect 5714 24360 6040 24378
rect 5714 24310 6015 24360
rect 6032 24310 6040 24360
rect 5714 24292 6040 24310
rect 5714 24218 6040 24236
rect 5714 24168 6015 24218
rect 6032 24168 6040 24218
rect 5714 24150 6040 24168
rect 5714 24076 6040 24094
rect 5714 24026 6015 24076
rect 6032 24026 6040 24076
rect 5714 24008 6040 24026
rect 5714 23934 6040 23952
rect 5714 23884 6015 23934
rect 6032 23884 6040 23934
rect 5714 23866 6040 23884
rect 5714 23792 6040 23810
rect 5714 23742 6015 23792
rect 6032 23742 6040 23792
rect 5714 23724 6040 23742
rect 5714 23650 6040 23668
rect 5714 23600 6015 23650
rect 6032 23600 6040 23650
rect 5714 23582 6040 23600
rect 5714 23508 6040 23526
rect 5714 23458 6015 23508
rect 6032 23458 6040 23508
rect 5714 23440 6040 23458
rect 5714 23366 6040 23384
rect 5714 23316 6015 23366
rect 6032 23316 6040 23366
rect 5714 23298 6040 23316
rect 5714 23224 6040 23242
rect 5714 23174 6015 23224
rect 6032 23174 6040 23224
rect 5714 23156 6040 23174
rect 5714 23082 6040 23100
rect 5714 23032 6015 23082
rect 6032 23032 6040 23082
rect 5714 23014 6040 23032
rect 5714 22940 6040 22958
rect 5714 22890 6015 22940
rect 6032 22890 6040 22940
rect 5714 22872 6040 22890
rect 5714 22798 6040 22816
rect 5714 22748 6015 22798
rect 6032 22748 6040 22798
rect 5714 22730 6040 22748
rect 5714 22656 6040 22674
rect 5714 22606 6015 22656
rect 6032 22606 6040 22656
rect 5714 22588 6040 22606
rect 5714 22514 6040 22532
rect 5714 22464 6015 22514
rect 6032 22464 6040 22514
rect 5714 22446 6040 22464
rect 5714 22372 6040 22390
rect 5714 22322 6015 22372
rect 6032 22322 6040 22372
rect 5714 22304 6040 22322
rect 5714 22230 6040 22248
rect 5714 22180 6015 22230
rect 6032 22180 6040 22230
rect 5714 22162 6040 22180
rect 5714 22088 6040 22106
rect 5714 22038 6015 22088
rect 6032 22038 6040 22088
rect 5714 22020 6040 22038
rect 5714 21946 6040 21964
rect 5714 21896 6015 21946
rect 6032 21896 6040 21946
rect 5714 21878 6040 21896
rect 5714 21804 6040 21822
rect 5714 21754 6015 21804
rect 6032 21754 6040 21804
rect 5714 21736 6040 21754
rect 5714 21662 6040 21680
rect 5714 21612 6015 21662
rect 6032 21612 6040 21662
rect 5714 21594 6040 21612
rect 5714 21520 6040 21538
rect 5714 21470 6015 21520
rect 6032 21470 6040 21520
rect 5714 21452 6040 21470
rect 5714 21378 6040 21396
rect 5714 21328 6015 21378
rect 6032 21328 6040 21378
rect 5714 21310 6040 21328
rect 5714 21236 6040 21254
rect 5714 21186 6015 21236
rect 6032 21186 6040 21236
rect 5714 21168 6040 21186
rect 5714 21094 6040 21112
rect 5714 21044 6015 21094
rect 6032 21044 6040 21094
rect 5714 21026 6040 21044
rect 5714 20952 6040 20970
rect 5714 20902 6015 20952
rect 6032 20902 6040 20952
rect 5714 20884 6040 20902
rect 5714 20810 6040 20828
rect 5714 20760 6015 20810
rect 6032 20760 6040 20810
rect 5714 20742 6040 20760
rect 5714 20668 6040 20686
rect 5714 20618 6015 20668
rect 6032 20618 6040 20668
rect 5714 20600 6040 20618
rect 5714 20526 6040 20544
rect 5714 20476 6015 20526
rect 6032 20476 6040 20526
rect 5714 20458 6040 20476
rect 5714 20384 6040 20402
rect 5714 20334 6015 20384
rect 6032 20334 6040 20384
rect 5714 20316 6040 20334
rect 5714 20242 6040 20260
rect 5714 20192 6015 20242
rect 6032 20192 6040 20242
rect 5714 20174 6040 20192
rect 5714 20100 6040 20118
rect 5714 20050 6015 20100
rect 6032 20050 6040 20100
rect 5714 20032 6040 20050
rect 5714 19958 6040 19976
rect 5714 19908 6015 19958
rect 6032 19908 6040 19958
rect 5714 19890 6040 19908
rect 5714 19816 6040 19834
rect 5714 19766 6015 19816
rect 6032 19766 6040 19816
rect 5714 19748 6040 19766
rect 5714 19674 6040 19692
rect 5714 19624 6015 19674
rect 6032 19624 6040 19674
rect 5714 19606 6040 19624
rect 5714 19532 6040 19550
rect 5714 19482 6015 19532
rect 6032 19482 6040 19532
rect 5714 19464 6040 19482
rect 5714 19390 6040 19408
rect 5714 19340 6015 19390
rect 6032 19340 6040 19390
rect 5714 19322 6040 19340
rect 5714 19248 6040 19266
rect 5714 19198 6015 19248
rect 6032 19198 6040 19248
rect 5714 19180 6040 19198
rect 5714 19106 6040 19124
rect 5714 19056 6015 19106
rect 6032 19056 6040 19106
rect 5714 19038 6040 19056
rect 5714 18964 6040 18982
rect 5714 18914 6015 18964
rect 6032 18914 6040 18964
rect 5714 18896 6040 18914
rect 5714 18822 6040 18840
rect 5714 18772 6015 18822
rect 6032 18772 6040 18822
rect 5714 18754 6040 18772
rect 5714 18680 6040 18698
rect 5714 18630 6015 18680
rect 6032 18630 6040 18680
rect 5714 18612 6040 18630
rect 5714 18538 6040 18556
rect 5714 18488 6015 18538
rect 6032 18488 6040 18538
rect 5714 18470 6040 18488
rect 5714 18396 6040 18414
rect 5714 18346 6015 18396
rect 6032 18346 6040 18396
rect 5714 18328 6040 18346
rect 5714 18254 6040 18272
rect 5714 18204 6015 18254
rect 6032 18204 6040 18254
rect 5714 18186 6040 18204
rect 5714 18112 6040 18130
rect 5714 18062 6015 18112
rect 6032 18062 6040 18112
rect 5714 18044 6040 18062
rect 5714 17970 6040 17988
rect 5714 17920 6015 17970
rect 6032 17920 6040 17970
rect 5714 17902 6040 17920
rect 5714 17828 6040 17846
rect 5714 17778 6015 17828
rect 6032 17778 6040 17828
rect 5714 17760 6040 17778
rect 5714 17686 6040 17704
rect 5714 17636 6015 17686
rect 6032 17636 6040 17686
rect 5714 17618 6040 17636
rect 5714 17544 6040 17562
rect 5714 17494 6015 17544
rect 6032 17494 6040 17544
rect 5714 17476 6040 17494
rect 5714 17402 6040 17420
rect 5714 17352 6015 17402
rect 6032 17352 6040 17402
rect 5714 17334 6040 17352
rect 5714 17260 6040 17278
rect 5714 17210 6015 17260
rect 6032 17210 6040 17260
rect 5714 17192 6040 17210
rect 5714 17118 6040 17136
rect 5714 17068 6015 17118
rect 6032 17068 6040 17118
rect 5714 17050 6040 17068
rect 5714 16976 6040 16994
rect 5714 16926 6015 16976
rect 6032 16926 6040 16976
rect 5714 16908 6040 16926
rect 5714 16834 6040 16852
rect 5714 16784 6015 16834
rect 6032 16784 6040 16834
rect 5714 16766 6040 16784
rect 5714 16692 6040 16710
rect 5714 16642 6015 16692
rect 6032 16642 6040 16692
rect 5714 16624 6040 16642
rect 5714 16550 6040 16568
rect 5714 16500 6015 16550
rect 6032 16500 6040 16550
rect 5714 16482 6040 16500
rect 5714 16408 6040 16426
rect 5714 16358 6015 16408
rect 6032 16358 6040 16408
rect 5714 16340 6040 16358
rect 5714 16266 6040 16284
rect 5714 16216 6015 16266
rect 6032 16216 6040 16266
rect 5714 16198 6040 16216
rect 5714 16124 6040 16142
rect 5714 16074 6015 16124
rect 6032 16074 6040 16124
rect 5714 16056 6040 16074
rect 5714 15982 6040 16000
rect 5714 15932 6015 15982
rect 6032 15932 6040 15982
rect 5714 15914 6040 15932
rect 5714 15840 6040 15858
rect 5714 15790 6015 15840
rect 6032 15790 6040 15840
rect 5714 15772 6040 15790
rect 5714 15698 6040 15716
rect 5714 15648 6015 15698
rect 6032 15648 6040 15698
rect 5714 15630 6040 15648
rect 5714 15556 6040 15574
rect 5714 15506 6015 15556
rect 6032 15506 6040 15556
rect 5714 15488 6040 15506
rect 5714 15414 6040 15432
rect 5714 15364 6015 15414
rect 6032 15364 6040 15414
rect 5714 15346 6040 15364
rect 5714 15272 6040 15290
rect 5714 15222 6015 15272
rect 6032 15222 6040 15272
rect 5714 15204 6040 15222
rect 5714 15130 6040 15148
rect 5714 15080 6015 15130
rect 6032 15080 6040 15130
rect 5714 15062 6040 15080
rect 5714 14988 6040 15006
rect 5714 14938 6015 14988
rect 6032 14938 6040 14988
rect 5714 14920 6040 14938
rect 5714 14846 6040 14864
rect 5714 14796 6015 14846
rect 6032 14796 6040 14846
rect 5714 14778 6040 14796
rect 5714 14704 6040 14722
rect 5714 14654 6015 14704
rect 6032 14654 6040 14704
rect 5714 14636 6040 14654
rect 5714 14562 6040 14580
rect 5714 14512 6015 14562
rect 6032 14512 6040 14562
rect 5714 14494 6040 14512
rect 5714 14420 6040 14438
rect 5714 14370 6015 14420
rect 6032 14370 6040 14420
rect 5714 14352 6040 14370
rect 5714 14278 6040 14296
rect 5714 14228 6015 14278
rect 6032 14228 6040 14278
rect 5714 14210 6040 14228
rect 5714 14136 6040 14154
rect 5714 14086 6015 14136
rect 6032 14086 6040 14136
rect 5714 14068 6040 14086
rect 5714 13994 6040 14012
rect 5714 13944 6015 13994
rect 6032 13944 6040 13994
rect 5714 13926 6040 13944
rect 5714 13852 6040 13870
rect 5714 13802 6015 13852
rect 6032 13802 6040 13852
rect 5714 13784 6040 13802
rect 5714 13710 6040 13728
rect 5714 13660 6015 13710
rect 6032 13660 6040 13710
rect 5714 13642 6040 13660
rect 5714 13568 6040 13586
rect 5714 13518 6015 13568
rect 6032 13518 6040 13568
rect 5714 13500 6040 13518
rect 5714 13426 6040 13444
rect 5714 13376 6015 13426
rect 6032 13376 6040 13426
rect 5714 13358 6040 13376
rect 5714 13284 6040 13302
rect 5714 13234 6015 13284
rect 6032 13234 6040 13284
rect 5714 13216 6040 13234
rect 5714 13142 6040 13160
rect 5714 13092 6015 13142
rect 6032 13092 6040 13142
rect 5714 13074 6040 13092
rect 5714 13000 6040 13018
rect 5714 12950 6015 13000
rect 6032 12950 6040 13000
rect 5714 12932 6040 12950
rect 5714 12858 6040 12876
rect 5714 12808 6015 12858
rect 6032 12808 6040 12858
rect 5714 12790 6040 12808
rect 5714 12716 6040 12734
rect 5714 12666 6015 12716
rect 6032 12666 6040 12716
rect 5714 12648 6040 12666
rect 5714 12574 6040 12592
rect 5714 12524 6015 12574
rect 6032 12524 6040 12574
rect 5714 12506 6040 12524
rect 5714 12432 6040 12450
rect 5714 12382 6015 12432
rect 6032 12382 6040 12432
rect 5714 12364 6040 12382
rect 5714 12290 6040 12308
rect 5714 12240 6015 12290
rect 6032 12240 6040 12290
rect 5714 12222 6040 12240
rect 5714 12148 6040 12166
rect 5714 12098 6015 12148
rect 6032 12098 6040 12148
rect 5714 12080 6040 12098
rect 5714 12006 6040 12024
rect 5714 11956 6015 12006
rect 6032 11956 6040 12006
rect 5714 11938 6040 11956
rect 5714 11864 6040 11882
rect 5714 11814 6015 11864
rect 6032 11814 6040 11864
rect 5714 11796 6040 11814
rect 5714 11722 6040 11740
rect 5714 11672 6015 11722
rect 6032 11672 6040 11722
rect 5714 11654 6040 11672
rect 5714 11580 6040 11598
rect 5714 11530 6015 11580
rect 6032 11530 6040 11580
rect 5714 11512 6040 11530
rect 5714 11438 6040 11456
rect 5714 11388 6015 11438
rect 6032 11388 6040 11438
rect 5714 11370 6040 11388
rect 5714 11296 6040 11314
rect 5714 11246 6015 11296
rect 6032 11246 6040 11296
rect 5714 11228 6040 11246
rect 5714 11154 6040 11172
rect 5714 11104 6015 11154
rect 6032 11104 6040 11154
rect 5714 11086 6040 11104
rect 5714 11012 6040 11030
rect 5714 10962 6015 11012
rect 6032 10962 6040 11012
rect 5714 10944 6040 10962
rect 5714 10870 6040 10888
rect 5714 10820 6015 10870
rect 6032 10820 6040 10870
rect 5714 10802 6040 10820
rect 5714 10728 6040 10746
rect 5714 10678 6015 10728
rect 6032 10678 6040 10728
rect 5714 10660 6040 10678
rect 5714 10586 6040 10604
rect 5714 10536 6015 10586
rect 6032 10536 6040 10586
rect 5714 10518 6040 10536
rect 5714 10444 6040 10462
rect 5714 10394 6015 10444
rect 6032 10394 6040 10444
rect 5714 10376 6040 10394
rect 5714 10302 6040 10320
rect 5714 10252 6015 10302
rect 6032 10252 6040 10302
rect 5714 10234 6040 10252
rect 5714 10160 6040 10178
rect 5714 10110 6015 10160
rect 6032 10110 6040 10160
rect 5714 10092 6040 10110
rect 5714 10018 6040 10036
rect 5714 9968 6015 10018
rect 6032 9968 6040 10018
rect 5714 9950 6040 9968
rect 5714 9876 6040 9894
rect 5714 9826 6015 9876
rect 6032 9826 6040 9876
rect 5714 9808 6040 9826
rect 5714 9734 6040 9752
rect 5714 9684 6015 9734
rect 6032 9684 6040 9734
rect 5714 9666 6040 9684
rect 5714 9592 6040 9610
rect 5714 9542 6015 9592
rect 6032 9542 6040 9592
rect 5714 9524 6040 9542
rect 5714 9450 6040 9468
rect 5714 9400 6015 9450
rect 6032 9400 6040 9450
rect 5714 9382 6040 9400
rect 5714 9308 6040 9326
rect 5714 9258 6015 9308
rect 6032 9258 6040 9308
rect 5714 9240 6040 9258
rect 5714 9166 6040 9184
rect 5714 9116 6015 9166
rect 6032 9116 6040 9166
rect 5714 9098 6040 9116
rect 5714 9024 6040 9042
rect 5714 8974 6015 9024
rect 6032 8974 6040 9024
rect 5714 8956 6040 8974
rect 5714 8882 6040 8900
rect 5714 8832 6015 8882
rect 6032 8832 6040 8882
rect 5714 8814 6040 8832
rect 5714 8740 6040 8758
rect 5714 8690 6015 8740
rect 6032 8690 6040 8740
rect 5714 8672 6040 8690
rect 5714 8598 6040 8616
rect 5714 8548 6015 8598
rect 6032 8548 6040 8598
rect 5714 8530 6040 8548
rect 5714 8456 6040 8474
rect 5714 8406 6015 8456
rect 6032 8406 6040 8456
rect 5714 8388 6040 8406
rect 5714 8314 6040 8332
rect 5714 8264 6015 8314
rect 6032 8264 6040 8314
rect 5714 8246 6040 8264
rect 5714 8172 6040 8190
rect 5714 8122 6015 8172
rect 6032 8122 6040 8172
rect 5714 8104 6040 8122
rect 5714 8030 6040 8048
rect 5714 7980 6015 8030
rect 6032 7980 6040 8030
rect 5714 7962 6040 7980
rect 5714 7888 6040 7906
rect 5714 7838 6015 7888
rect 6032 7838 6040 7888
rect 5714 7820 6040 7838
rect 5714 7746 6040 7764
rect 5714 7696 6015 7746
rect 6032 7696 6040 7746
rect 5714 7678 6040 7696
rect 5714 7604 6040 7622
rect 5714 7554 6015 7604
rect 6032 7554 6040 7604
rect 5714 7536 6040 7554
rect 5714 7462 6040 7480
rect 5714 7412 6015 7462
rect 6032 7412 6040 7462
rect 5714 7394 6040 7412
rect 5714 7320 6040 7338
rect 5714 7270 6015 7320
rect 6032 7270 6040 7320
rect 5714 7252 6040 7270
rect 5714 7178 6040 7196
rect 5714 7128 6015 7178
rect 6032 7128 6040 7178
rect 5714 7110 6040 7128
rect 5714 7036 6040 7054
rect 5714 6986 6015 7036
rect 6032 6986 6040 7036
rect 5714 6968 6040 6986
rect 5714 6894 6040 6912
rect 5714 6844 6015 6894
rect 6032 6844 6040 6894
rect 5714 6826 6040 6844
rect 5714 6752 6040 6770
rect 5714 6702 6015 6752
rect 6032 6702 6040 6752
rect 5714 6684 6040 6702
rect 5714 6610 6040 6628
rect 5714 6560 6015 6610
rect 6032 6560 6040 6610
rect 5714 6542 6040 6560
rect 5714 6468 6040 6486
rect 5714 6418 6015 6468
rect 6032 6418 6040 6468
rect 5714 6400 6040 6418
rect 5714 6326 6040 6344
rect 5714 6276 6015 6326
rect 6032 6276 6040 6326
rect 5714 6258 6040 6276
rect 5714 6184 6040 6202
rect 5714 6134 6015 6184
rect 6032 6134 6040 6184
rect 5714 6116 6040 6134
rect 5714 6042 6040 6060
rect 5714 5992 6015 6042
rect 6032 5992 6040 6042
rect 5714 5974 6040 5992
rect 5714 5900 6040 5918
rect 5714 5850 6015 5900
rect 6032 5850 6040 5900
rect 5714 5832 6040 5850
rect 5714 5758 6040 5776
rect 5714 5708 6015 5758
rect 6032 5708 6040 5758
rect 5714 5690 6040 5708
rect 5714 5616 6040 5634
rect 5714 5566 6015 5616
rect 6032 5566 6040 5616
rect 5714 5548 6040 5566
rect 5714 5474 6040 5492
rect 5714 5424 6015 5474
rect 6032 5424 6040 5474
rect 5714 5406 6040 5424
rect 5714 5332 6040 5350
rect 5714 5282 6015 5332
rect 6032 5282 6040 5332
rect 5714 5264 6040 5282
rect 5714 5190 6040 5208
rect 5714 5140 6015 5190
rect 6032 5140 6040 5190
rect 5714 5122 6040 5140
rect 5714 5048 6040 5066
rect 5714 4998 6015 5048
rect 6032 4998 6040 5048
rect 5714 4980 6040 4998
rect 5714 4906 6040 4924
rect 5714 4856 6015 4906
rect 6032 4856 6040 4906
rect 5714 4838 6040 4856
rect 5714 4764 6040 4782
rect 5714 4714 6015 4764
rect 6032 4714 6040 4764
rect 5714 4696 6040 4714
rect 5714 4622 6040 4640
rect 5714 4572 6015 4622
rect 6032 4572 6040 4622
rect 5714 4554 6040 4572
rect 5714 4480 6040 4498
rect 5714 4430 6015 4480
rect 6032 4430 6040 4480
rect 5714 4412 6040 4430
rect 5714 4338 6040 4356
rect 5714 4288 6015 4338
rect 6032 4288 6040 4338
rect 5714 4270 6040 4288
rect 5714 4196 6040 4214
rect 5714 4146 6015 4196
rect 6032 4146 6040 4196
rect 5714 4128 6040 4146
rect 5714 4054 6040 4072
rect 5714 4004 6015 4054
rect 6032 4004 6040 4054
rect 5714 3986 6040 4004
rect 5714 3912 6040 3930
rect 5714 3862 6015 3912
rect 6032 3862 6040 3912
rect 5714 3844 6040 3862
rect 5714 3770 6040 3788
rect 5714 3720 6015 3770
rect 6032 3720 6040 3770
rect 5714 3702 6040 3720
rect 5714 3628 6040 3646
rect 5714 3578 6015 3628
rect 6032 3578 6040 3628
rect 5714 3560 6040 3578
rect 5714 3486 6040 3504
rect 5714 3436 6015 3486
rect 6032 3436 6040 3486
rect 5714 3418 6040 3436
rect 5714 3344 6040 3362
rect 5714 3294 6015 3344
rect 6032 3294 6040 3344
rect 5714 3276 6040 3294
rect 5714 3202 6040 3220
rect 5714 3152 6015 3202
rect 6032 3152 6040 3202
rect 5714 3134 6040 3152
rect 5714 3060 6040 3078
rect 5714 3010 6015 3060
rect 6032 3010 6040 3060
rect 5714 2992 6040 3010
rect 5714 2918 6040 2936
rect 5714 2868 6015 2918
rect 6032 2868 6040 2918
rect 5714 2850 6040 2868
rect 5714 2776 6040 2794
rect 5714 2726 6015 2776
rect 6032 2726 6040 2776
rect 5714 2708 6040 2726
rect 5714 2634 6040 2652
rect 5714 2584 6015 2634
rect 6032 2584 6040 2634
rect 5714 2566 6040 2584
rect 5714 2492 6040 2510
rect 5714 2442 6015 2492
rect 6032 2442 6040 2492
rect 5714 2424 6040 2442
rect 5714 2350 6040 2368
rect 5714 2300 6015 2350
rect 6032 2300 6040 2350
rect 5714 2282 6040 2300
rect 5714 2208 6040 2226
rect 5714 2158 6015 2208
rect 6032 2158 6040 2208
rect 5714 2140 6040 2158
rect 5714 2066 6040 2084
rect 5714 2016 6015 2066
rect 6032 2016 6040 2066
rect 5714 1998 6040 2016
rect 5714 1924 6040 1942
rect 5714 1874 6015 1924
rect 6032 1874 6040 1924
rect 5714 1856 6040 1874
rect 5714 1782 6040 1800
rect 5714 1732 6015 1782
rect 6032 1732 6040 1782
rect 5714 1714 6040 1732
rect 5714 1640 6040 1658
rect 5714 1590 6015 1640
rect 6032 1590 6040 1640
rect 5714 1572 6040 1590
rect 5714 1498 6040 1516
rect 5714 1448 6015 1498
rect 6032 1448 6040 1498
rect 5714 1430 6040 1448
rect 5714 1356 6040 1374
rect 5714 1306 6015 1356
rect 6032 1306 6040 1356
rect 5714 1288 6040 1306
rect 5714 1214 6040 1232
rect 5714 1164 6015 1214
rect 6032 1164 6040 1214
rect 5714 1146 6040 1164
rect 5714 1072 6040 1090
rect 5714 1022 6015 1072
rect 6032 1022 6040 1072
rect 5714 1004 6040 1022
rect 5714 930 6040 948
rect 5714 880 6015 930
rect 6032 880 6040 930
rect 5714 862 6040 880
rect 5714 788 6040 806
rect 5714 738 6015 788
rect 6032 738 6040 788
rect 5714 720 6040 738
rect 5714 646 6040 664
rect 5714 596 6015 646
rect 6032 596 6040 646
rect 5714 578 6040 596
rect 5714 504 6040 522
rect 5714 454 6015 504
rect 6032 454 6040 504
rect 5714 436 6040 454
rect 5714 362 6040 380
rect 5714 312 6015 362
rect 6032 312 6040 362
rect 5714 294 6040 312
rect 5714 220 6040 238
rect 5714 170 6015 220
rect 6032 170 6040 220
rect 5714 152 6040 170
rect 6088 80 6196 92
rect 6088 60 6198 80
rect 6088 6 6108 60
rect 6174 6 6198 60
rect 6088 -2 6198 6
rect 6428 75 6536 94
rect 6428 9 6440 75
rect 6506 9 6536 75
rect 6428 0 6536 9
rect 6592 73 6700 96
rect 6592 7 6606 73
rect 6672 7 6700 73
rect 6592 2 6700 7
rect 6920 67 7028 100
rect 6920 13 6938 67
rect 7004 13 7028 67
rect 6920 6 7028 13
rect 7090 66 7198 94
rect 7418 72 7526 92
rect 7090 60 7210 66
rect 7090 6 7104 60
rect 7170 6 7210 60
rect 6600 1 6678 2
rect 50 -78 106 -72
rect 5548 -78 5604 -66
rect 50 -84 5554 -78
rect 50 -128 56 -84
rect 100 -128 5554 -84
rect 50 -134 5554 -128
rect 5598 -134 5604 -78
rect 50 -140 106 -134
rect 5548 -146 5604 -134
rect 6108 -205 6174 -2
rect 5727 -271 6174 -205
rect 5727 -659 5793 -271
rect 6440 -311 6506 0
rect 5727 -713 5733 -659
rect 5787 -713 5793 -659
rect 5727 -725 5793 -713
rect 6033 -377 6506 -311
rect 6033 -661 6099 -377
rect 6606 -439 6672 1
rect 6033 -715 6039 -661
rect 6093 -715 6099 -661
rect 6033 -727 6099 -715
rect 6335 -505 6672 -439
rect 6335 -661 6401 -505
rect 6938 -523 7004 6
rect 7090 0 7210 6
rect 6829 -589 7004 -523
rect 7141 -466 7210 0
rect 7418 6 7436 72
rect 7502 6 7526 72
rect 7418 -2 7526 6
rect 7586 60 7694 94
rect 7930 81 8038 90
rect 7928 75 8038 81
rect 7586 6 7602 60
rect 7668 6 7694 60
rect 7586 0 7694 6
rect 7877 9 7934 75
rect 8000 9 8038 75
rect 6829 -653 6895 -589
rect 6335 -715 6341 -661
rect 6395 -715 6401 -661
rect 6335 -727 6401 -715
rect 6641 -659 6895 -653
rect 7141 -657 7207 -466
rect 6641 -713 6653 -659
rect 6707 -713 6895 -659
rect 6641 -719 6895 -713
rect 6955 -663 7207 -657
rect 7436 -663 7502 -2
rect 7602 -655 7668 0
rect 6955 -717 6967 -663
rect 7021 -717 7207 -663
rect 6955 -723 7207 -717
rect 7251 -669 7502 -663
rect 7251 -723 7263 -669
rect 7317 -723 7502 -669
rect 7553 -661 7668 -655
rect 7553 -715 7565 -661
rect 7619 -715 7668 -661
rect 7553 -721 7668 -715
rect 7877 -4 8038 9
rect 7877 -661 7943 -4
rect 7877 -715 7883 -661
rect 7937 -715 7943 -661
rect 7251 -729 7502 -723
rect 7877 -727 7943 -715
<< via1 >>
rect -222 145220 -164 145276
rect -161 142319 -95 142385
rect -177 139064 -111 139130
rect -138 135867 -86 135919
rect -135 132593 -69 132659
rect -119 129359 -53 129425
rect -139 126117 -73 126183
rect -157 122885 -91 122951
rect -524 119528 -446 119534
rect -524 119462 -518 119528
rect -518 119462 -452 119528
rect -452 119462 -446 119528
rect -524 119456 -446 119462
rect -637 118821 -571 118827
rect -637 118767 -631 118821
rect -631 118767 -577 118821
rect -577 118767 -571 118821
rect -637 118761 -571 118767
rect -619 118419 -553 118425
rect -619 118365 -613 118419
rect -613 118365 -559 118419
rect -559 118365 -553 118419
rect -619 118359 -553 118365
rect -637 118185 -571 118191
rect -637 118131 -631 118185
rect -631 118131 -577 118185
rect -577 118131 -571 118185
rect -637 118125 -571 118131
rect -627 117805 -545 117811
rect -627 117735 -621 117805
rect -621 117735 -551 117805
rect -551 117735 -545 117805
rect -627 117729 -545 117735
rect -477 117370 -411 117376
rect -477 117316 -471 117370
rect -471 117316 -417 117370
rect -417 117316 -411 117370
rect -477 117310 -411 117316
rect -398 114316 -346 114390
rect -401 111057 -335 111123
rect -394 107814 -338 107894
<< metal2 >>
rect 436 146748 502 146814
rect 700 146654 766 146720
rect 957 146626 1023 146635
rect 957 146560 1030 146626
rect 957 145622 1023 146560
rect 1222 146532 1289 146535
rect 1222 146466 1294 146532
rect 953 145566 962 145622
rect 1018 145566 1027 145622
rect 957 145561 1023 145566
rect -232 145276 -152 145286
rect -232 145220 -222 145276
rect -164 145220 -152 145276
rect -232 145210 -152 145220
rect -172 142385 -86 142396
rect -172 142319 -161 142385
rect -95 142319 -86 142385
rect 1222 142381 1289 146466
rect 1479 146436 1550 146442
rect 1479 146370 1562 146436
rect 1216 142324 1225 142381
rect 1286 142324 1295 142381
rect 1222 142319 1289 142324
rect -172 142310 -86 142319
rect -182 139130 -104 139138
rect -182 139064 -177 139130
rect -111 139064 -104 139130
rect -182 139058 -104 139064
rect 1479 139125 1550 146370
rect 1756 146341 1822 146344
rect 1479 139069 1486 139125
rect 1542 139069 1550 139125
rect 1479 139050 1550 139069
rect 1753 146278 1822 146341
rect -150 135921 -74 135932
rect -150 135865 -140 135921
rect -84 135865 -74 135921
rect -150 135856 -74 135865
rect 1753 135921 1819 146278
rect 1753 135865 1758 135921
rect 1814 135865 1819 135921
rect 1753 135860 1819 135865
rect 1758 135856 1814 135860
rect -144 132659 -60 132668
rect -144 132593 -135 132659
rect -69 132593 -60 132659
rect -144 132582 -60 132593
rect 2020 132649 2086 146250
rect 2020 132584 2086 132593
rect 2284 131159 2350 146156
rect 2279 131099 2350 131159
rect 2554 131145 2621 146069
rect 2819 145902 2893 145958
rect -128 129425 -44 129434
rect -128 129359 -119 129425
rect -53 129359 -44 129425
rect 2279 129420 2345 131099
rect 2279 129364 2284 129420
rect 2340 129364 2345 129420
rect 2279 129359 2345 129364
rect 2533 131049 2621 131145
rect -128 129350 -44 129359
rect 2284 129355 2340 129359
rect -144 126183 -60 126192
rect -144 126117 -139 126183
rect -73 126117 -60 126183
rect -144 126108 -60 126117
rect 2533 126173 2599 131049
rect 2837 130831 2893 145902
rect 2533 126117 2538 126173
rect 2594 126117 2599 126173
rect 2533 126112 2599 126117
rect 2538 126108 2594 126112
rect -166 122951 -82 122960
rect -166 122885 -157 122951
rect -91 122885 -82 122951
rect 2829 122946 2895 130831
rect 2829 122890 2834 122946
rect 2890 122890 2895 122946
rect 2829 122885 2895 122890
rect -166 122876 -82 122885
rect 2834 122881 2890 122885
rect -397 120191 -331 120301
rect -518 120125 -331 120191
rect -518 119540 -452 120125
rect -532 119534 -438 119540
rect -532 119456 -524 119534
rect -446 119456 -438 119534
rect -532 119450 -438 119456
rect -643 118761 -637 118827
rect -571 118761 -289 118827
rect -626 118425 -546 118432
rect -626 118359 -619 118425
rect -553 118359 -546 118425
rect -626 118352 -546 118359
rect -644 118191 -564 118198
rect -644 118125 -637 118191
rect -571 118125 -564 118191
rect -644 118118 -564 118125
rect -634 117811 -538 117818
rect -634 117729 -627 117811
rect -545 117729 -538 117811
rect -634 117722 -538 117729
rect -355 117376 -289 118761
rect -483 117310 -477 117376
rect -411 117310 -289 117376
rect -414 114390 -336 114400
rect -414 114316 -402 114390
rect -346 114316 -336 114390
rect -414 114302 -336 114316
rect -410 111123 -330 111132
rect -410 111057 -401 111123
rect -335 111057 -330 111123
rect -410 111048 -330 111057
rect -406 107894 -332 107904
rect -406 107814 -394 107894
rect -338 107814 -332 107894
rect -406 107802 -332 107814
rect -398 105166 -334 105238
<< via2 >>
rect 962 145566 1018 145622
rect -222 145220 -164 145276
rect -161 142319 -95 142385
rect 1225 142324 1286 142381
rect -172 139069 -116 139125
rect 1486 139069 1542 139125
rect -140 135919 -84 135921
rect -140 135867 -138 135919
rect -138 135867 -86 135919
rect -86 135867 -84 135919
rect -140 135865 -84 135867
rect 1758 135865 1814 135921
rect -135 132593 -69 132659
rect 2020 132593 2086 132649
rect -119 129359 -53 129425
rect 2284 129364 2340 129420
rect -139 126117 -73 126173
rect 2538 126117 2594 126173
rect -157 122885 -91 122951
rect 2834 122890 2890 122946
rect -614 118364 -558 118420
rect -632 118130 -576 118186
rect -622 117734 -550 117806
rect -402 114316 -398 114390
rect -398 114316 -346 114390
rect -401 111057 -335 111123
rect -394 107814 -338 107894
<< metal3 >>
rect -50 145622 1028 145627
rect -50 145566 962 145622
rect 1018 145566 1028 145622
rect -50 145561 1028 145566
rect -232 145281 -152 145286
rect -49 145281 17 145561
rect -232 145276 17 145281
rect -232 145220 -222 145276
rect -164 145220 17 145276
rect -232 145215 17 145220
rect -232 145210 -152 145215
rect -166 142385 -90 142390
rect 851 142385 1292 142386
rect -166 142319 -161 142385
rect -95 142381 1292 142385
rect -95 142324 1225 142381
rect 1286 142324 1292 142381
rect -95 142319 1292 142324
rect -166 142314 -90 142319
rect -181 139125 1547 139130
rect -181 139069 -172 139125
rect -116 139069 1486 139125
rect 1542 139069 1547 139125
rect -181 139064 1547 139069
rect -145 135923 -79 135926
rect 1477 135923 1819 135926
rect -145 135921 1819 135923
rect -145 135865 -140 135921
rect -84 135865 1758 135921
rect 1814 135865 1819 135921
rect -145 135863 1819 135865
rect -145 135860 -79 135863
rect 1477 135860 1819 135863
rect -140 132659 -64 132664
rect -140 132593 -135 132659
rect -69 132654 803 132659
rect -69 132649 2091 132654
rect -69 132593 2020 132649
rect 2086 132593 2091 132649
rect -140 132588 -64 132593
rect 621 132588 2091 132593
rect -124 129425 -48 129430
rect -124 129359 -119 129425
rect -53 129420 2345 129425
rect -53 129364 2284 129420
rect 2340 129364 2345 129420
rect -53 129359 2345 129364
rect -124 129354 -48 129359
rect -144 126173 2599 126178
rect -144 126117 -139 126173
rect -73 126117 2538 126173
rect 2594 126117 2599 126173
rect -144 126112 2599 126117
rect -162 122951 -86 122956
rect -162 122885 -157 122951
rect -91 122946 2895 122951
rect -91 122890 2834 122946
rect 2890 122890 2895 122946
rect -91 122885 2895 122890
rect -162 122880 -86 122885
rect -540 118425 -335 118431
rect -619 118420 -335 118425
rect -619 118364 -614 118420
rect -558 118365 -335 118420
rect -558 118364 -540 118365
rect -619 118359 -540 118364
rect -881 118186 -571 118191
rect -881 118130 -632 118186
rect -576 118130 -571 118186
rect -881 118125 -571 118130
rect -881 111123 -815 118125
rect -717 117806 -545 117811
rect -717 117734 -622 117806
rect -550 117734 -545 117806
rect -717 117729 -545 117734
rect -717 111406 -635 117729
rect -401 114400 -335 118365
rect -414 114390 -335 114400
rect -414 114316 -402 114390
rect -346 114374 -335 114390
rect -346 114316 -336 114374
rect -414 114302 -336 114316
rect -722 111326 -716 111406
rect -636 111326 -630 111406
rect -717 111325 -635 111326
rect -406 111123 -330 111128
rect -881 111057 -401 111123
rect -335 111057 -330 111123
rect -406 111052 -330 111057
rect -717 110855 -635 110861
rect -717 107895 -635 110775
rect -406 107900 -332 107904
rect -410 107895 -328 107900
rect -717 107894 -328 107895
rect -717 107814 -394 107894
rect -338 107814 -328 107894
rect -717 107813 -328 107814
rect -410 107802 -328 107813
<< via3 >>
rect -716 111326 -636 111406
rect -717 110775 -635 110855
<< metal4 >>
rect -717 111406 -635 111407
rect -717 111326 -716 111406
rect -636 111326 -635 111406
rect -717 110856 -635 111326
rect -718 110855 -634 110856
rect -718 110775 -717 110855
rect -635 110775 -634 110855
rect -718 110774 -634 110775
use counter_4  counter_4_0
timestamp 1745485683
transform 0 -1 -40 1 0 105408
box -318 0 12226 976
use counter_8  counter_8_0
timestamp 1745486774
transform 0 -1 -40 1 0 120476
box -318 0 25180 976
use decoder_8  decoder_8_0
timestamp 1745492145
transform 1 0 238 0 1 145618
box -238 -145618 5702 1196
use inv  inv_0 ~/magic/library/mag
timestamp 1738780557
transform 0 -1 -40 1 0 119536
box -4 0 322 976
use inv  inv_1
timestamp 1738780557
transform 0 -1 -40 1 0 119844
box -4 0 322 976
use inv  inv_2
timestamp 1738780557
transform 1 0 6572 0 1 -1020
box -4 0 322 976
use inv  inv_3
timestamp 1738780557
transform 1 0 6264 0 1 -1020
box -4 0 322 976
use inv  inv_4
timestamp 1738780557
transform 1 0 7188 0 1 -1020
box -4 0 322 976
use inv  inv_5
timestamp 1738780557
transform 1 0 6880 0 1 -1020
box -4 0 322 976
use inv  inv_6
timestamp 1738780557
transform 1 0 5648 0 1 -1020
box -4 0 322 976
use inv  inv_7
timestamp 1738780557
transform 1 0 5956 0 1 -1020
box -4 0 322 976
use inv  inv_8
timestamp 1738780557
transform 1 0 7804 0 1 -1020
box -4 0 322 976
use inv  inv_9
timestamp 1738780557
transform 1 0 7496 0 1 -1020
box -4 0 322 976
use memory_8  memory_8_0
timestamp 1744679307
transform 1 0 6108 0 1 145480
box -134 -145474 1992 600
use mux4  mux4_0
timestamp 1745483395
transform 0 -1 -40 1 0 117626
box 0 0 1914 976
<< labels >>
flabel metal1 -202 119384 -137 119506 0 FreeSerif 160 270 0 0 Freq1
port 3 nsew
flabel metal2 -398 105166 -334 105238 0 FreeSerif 160 270 0 0 CLK
port 1 nsew
flabel metal1 -963 119428 -898 119550 0 FreeSerif 160 270 0 0 Freq0
port 2 nsew
flabel metal2 436 146748 502 146814 0 FreeSerif 160 0 0 0 Wave1
port 21 nsew
flabel metal2 700 146654 766 146720 0 FreeSerif 160 0 0 0 Wave0
port 20 nsew
flabel locali 5828 -674 5894 -472 0 FreeSerif 160 0 0 0 Y7
port 19 nsew
flabel locali 6136 -674 6202 -472 0 FreeSerif 160 0 0 0 Y6
port 18 nsew
flabel locali 6444 -674 6510 -472 0 FreeSerif 160 0 0 0 Y5
port 17 nsew
flabel locali 6752 -564 6818 -362 0 FreeSerif 160 0 0 0 Y4
port 16 nsew
flabel locali 7060 -584 7126 -382 0 FreeSerif 160 0 0 0 Y3
port 15 nsew
flabel locali 7368 -592 7434 -390 0 FreeSerif 160 0 0 0 Y2
port 14 nsew
flabel locali 7676 -594 7742 -392 0 FreeSerif 160 0 0 0 Y1
port 13 nsew
flabel locali 7984 -598 8050 -396 0 FreeSerif 160 0 0 0 Y0
port 12 nsew
<< end >>
