* NGSPICE file created from decoder_out.ext - technology: sky130A

*.subckt decoder_out A0 A1 A2 A3 word0 word1 word2 word3 word4 word5 word6 word7 word8
+ word9 word10 word11 word12 word13 word14 word15 VDD GND
X0 GND A0 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1 a_446_n626# A2 a_182_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2 a_50_n2046# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3 a_2292_n2330# a_2236_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4 GND A3 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5 word2 a_1708_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6 GND A0 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7 GND A2 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8 word14 A0 a_578_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9 a_446_n1478# A2 a_50_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10 GND A0 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11 a_182_n200# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12 a_314_n768# a_264_n66# a_182_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13 a_50_n2330# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14 GND A3 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15 a_1500_n1762# a_1444_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16 a_710_n1336# A1 a_446_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17 a_314_n1194# a_264_n66# a_182_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18 word7 a_792_n66# a_578_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19 GND A1 a_528_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X20 word7 a_1972_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X21 a_1708_164# A1 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X22 a_446_n484# A2 a_182_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X23 a_2292_n2188# a_2236_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X24 GND A3 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X25 a_578_n2330# a_528_n66# a_314_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X26 VDD A1 a_528_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X27 word9 a_792_n66# a_710_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X28 a_1708_164# A1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X29 a_50_n2188# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X30 GND A3 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X31 word0 A0 a_710_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X32 word13 a_1444_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X33 GND A1 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X34 word1 a_1444_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X35 GND A3 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X36 a_578_n2188# a_528_n66# a_314_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X37 a_710_n1478# A1 a_446_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X38 a_1500_n2330# a_1444_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X39 a_1500_n626# a_1444_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X40 GND A2 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X41 a_182_n342# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X42 word6 A0 a_578_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X43 word5 a_1444_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X44 GND A2 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X45 GND A2 a_264_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X46 a_182_n626# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X47 GND A1 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X48 word8 A0 a_710_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X49 VDD A2 a_264_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X50 word11 a_1708_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X51 GND A1 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X52 a_182_n910# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X53 a_578_n626# a_528_n66# a_446_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X54 word10 A0 a_578_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X55 a_314_n1904# a_264_n66# a_50_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X56 GND A2 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X57 a_2292_n1336# a_2236_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X58 a_2028_n1904# a_1972_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X59 a_446_n1762# A2 a_50_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X60 GND A0 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X61 a_182_n484# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X62 GND A2 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X63 a_50_n1336# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X64 a_2292_n1620# a_2236_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X65 a_578_n1052# a_528_n66# a_314_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X66 a_182_n768# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X67 a_710_n1904# A1 a_314_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X68 a_578_n484# a_528_n66# a_446_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X69 a_710_n200# A1 a_446_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X70 a_1764_n2330# a_1708_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X71 GND A2 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X72 word11 a_792_n66# a_578_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X73 a_50_n1620# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X74 a_2236_164# A3 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X75 word2 A0 a_578_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X76 a_1444_164# A0 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X77 a_2236_164# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X78 a_2292_n1478# a_2236_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X79 a_578_n1620# a_528_n66# a_446_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X80 GND A1 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X81 a_1444_164# A0 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X82 a_1764_n2188# a_1708_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X83 GND A1 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X84 GND A2 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X85 a_314_n2046# a_264_n66# a_50_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X86 word4 A0 a_710_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X87 word13 a_792_n66# a_710_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X88 a_50_n1478# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X89 a_2028_n2046# a_1972_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X90 a_578_n1194# a_528_n66# a_314_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X91 a_182_n1052# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X92 a_314_n2330# a_264_n66# a_50_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X93 word15 a_792_n66# a_578_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X94 GND A1 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X95 a_2028_n2330# a_1972_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X96 GND A0 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X97 a_710_n2046# A1 a_314_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X98 a_710_n342# A1 a_446_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X99 GND A0 a_792_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X100 word5 a_1972_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X101 a_1500_n1194# a_1444_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X102 VDD A0 a_792_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X103 word12 A0 a_710_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X104 a_314_n2188# a_264_n66# a_50_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X105 a_2028_n2188# a_1972_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X106 word9 a_1444_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X107 GND A1 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X108 GND A0 word14 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X109 a_182_n1194# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X110 GND A1 word13 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X111 a_710_n910# A1 a_314_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X112 a_446_n200# A2 a_182_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X113 word1 a_792_n66# a_710_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X114 GND A3 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X115 word4 a_1972_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X116 a_2292_n1904# a_2236_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X117 a_1764_n1052# a_1708_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X118 word3 a_792_n66# a_578_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X119 GND A3 a_0_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X120 GND A3 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X121 a_50_n1904# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X122 VDD A3 a_0_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X123 word5 a_792_n66# a_710_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X124 a_710_n768# A1 a_314_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X125 a_2292_n1762# a_2236_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X126 word10 a_1708_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X127 GND A2 word11 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X128 GND A3 word7 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X129 a_446_n1336# A2 a_50_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X130 a_50_n1762# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X131 a_314_n1052# a_264_n66# a_182_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X132 a_1764_n1194# a_1708_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X133 word3 a_1708_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X134 a_1972_164# A2 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X135 word6 a_1972_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X136 a_446_n1620# A2 a_50_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X137 GND A0 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X138 a_446_n342# A2 a_182_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X139 a_314_n910# a_264_n66# a_182_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X140 a_578_n1762# a_528_n66# a_446_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X141 a_2292_n2046# a_2236_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X142 a_1972_164# A2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X143 GND A0 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
*.ends

