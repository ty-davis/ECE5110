magic
tech sky130A
magscale 1 2
timestamp 1745486774
<< psubdiff >>
rect 22662 20 22682 76
<< locali >>
rect -314 864 22674 960
rect 22676 864 25180 960
rect 2685 693 2739 747
rect 5923 693 5977 747
rect 9161 693 9215 747
rect 12399 693 12453 747
rect 15637 693 15691 747
rect 18875 693 18929 747
rect 22113 693 22167 747
rect 3104 498 3170 692
rect 1010 374 1062 426
rect 4248 374 4300 426
rect 6342 474 6408 668
rect 9580 488 9646 682
rect 7486 374 7538 426
rect 10724 374 10776 426
rect 12818 474 12884 668
rect 16056 488 16122 682
rect 13962 374 14014 426
rect 17200 374 17252 426
rect 19294 474 19360 668
rect 22532 488 22598 682
rect 20438 374 20490 426
rect 23678 374 23730 426
rect 24856 370 24922 436
rect 1738 306 1792 358
rect 2788 304 3068 368
rect 3104 295 3343 361
rect 4976 306 5030 358
rect 6026 304 6306 368
rect 6342 291 6593 357
rect 8214 306 8268 358
rect 9264 304 9544 368
rect 9722 359 9819 361
rect 9580 295 9819 359
rect 11452 306 11506 358
rect 12502 304 12782 368
rect 9580 293 9722 295
rect 12818 291 13069 357
rect 14690 306 14744 358
rect 15740 304 16020 368
rect 16198 359 16295 361
rect 16056 295 16295 359
rect 17928 306 17982 358
rect 18978 304 19258 368
rect 16056 293 16198 295
rect 19294 291 19545 357
rect 21166 306 21220 358
rect 22216 304 22496 368
rect 22654 359 22696 360
rect 22532 293 22801 359
rect 24406 306 24460 358
rect 22654 292 22696 293
rect -314 0 25180 96
<< viali >>
rect 88 625 142 679
rect -130 414 -90 454
rect 2689 423 2743 477
rect 2202 384 2240 422
rect 5929 423 5983 477
rect 9165 427 9219 481
rect 5440 384 5478 422
rect 8678 384 8716 422
rect 12405 423 12459 477
rect 15641 427 15695 481
rect 11916 384 11954 422
rect 15154 384 15192 422
rect 18881 423 18935 477
rect 22117 427 22171 481
rect 18392 384 18430 422
rect 21630 384 21668 422
rect -231 299 -177 353
rect 2581 301 2635 355
rect 5819 301 5873 355
rect 9057 301 9111 355
rect 12295 301 12349 355
rect 15533 301 15587 355
rect 18771 301 18825 355
rect 22009 301 22063 355
<< metal1 >>
rect 82 679 148 691
rect 82 625 88 679
rect 142 625 148 679
rect 82 529 148 625
rect 407 531 413 597
rect 479 531 485 597
rect 2549 523 2555 589
rect 2621 523 2627 589
rect 3645 531 3651 597
rect 3717 531 3723 597
rect 2555 483 2621 523
rect 5804 521 5810 587
rect 5876 521 5882 587
rect 6883 531 6889 597
rect 6955 531 6961 597
rect 9040 521 9046 587
rect 9112 521 9118 587
rect 10121 531 10127 597
rect 10193 531 10199 597
rect 12280 521 12286 587
rect 12352 521 12358 587
rect 13359 531 13365 597
rect 13431 531 13437 597
rect 15516 521 15522 587
rect 15588 521 15594 587
rect 16597 531 16603 597
rect 16669 531 16675 597
rect 18756 521 18762 587
rect 18828 521 18834 587
rect 19835 531 19841 597
rect 19907 531 19913 597
rect 21992 521 21998 587
rect 22064 521 22070 587
rect 23075 531 23153 597
rect 5810 483 5876 521
rect 9046 487 9112 521
rect 2555 477 2755 483
rect -136 460 -84 466
rect -136 402 -84 408
rect 2188 422 2457 436
rect 2188 384 2202 422
rect 2240 384 2457 422
rect 2555 423 2689 477
rect 2743 423 2755 477
rect 5810 477 5995 483
rect 2555 417 2755 423
rect 2188 370 2457 384
rect 5426 422 5695 436
rect 5426 384 5440 422
rect 5478 384 5695 422
rect 5810 423 5929 477
rect 5983 423 5995 477
rect 9046 481 9231 487
rect 5810 417 5995 423
rect 5426 370 5695 384
rect 8664 422 8933 436
rect 8664 384 8678 422
rect 8716 384 8933 422
rect 9046 427 9165 481
rect 9219 427 9231 481
rect 12286 483 12352 521
rect 15522 487 15588 521
rect 12286 477 12471 483
rect 9046 421 9231 427
rect 8664 370 8933 384
rect 11902 422 12171 436
rect 11902 384 11916 422
rect 11954 384 12171 422
rect 12286 423 12405 477
rect 12459 423 12471 477
rect 15522 481 15707 487
rect 12286 417 12471 423
rect 11902 370 12171 384
rect 15140 422 15409 436
rect 15140 384 15154 422
rect 15192 384 15409 422
rect 15522 427 15641 481
rect 15695 427 15707 481
rect 18762 483 18828 521
rect 21998 487 22064 521
rect 18762 477 18947 483
rect 15522 421 15707 427
rect 15140 370 15409 384
rect 18378 422 18647 436
rect 18378 384 18392 422
rect 18430 384 18647 422
rect 18762 423 18881 477
rect 18935 423 18947 477
rect 21998 481 22183 487
rect 18762 417 18947 423
rect 18378 370 18647 384
rect 21616 422 21885 436
rect 21616 384 21630 422
rect 21668 384 21885 422
rect 21998 427 22117 481
rect 22171 427 22183 481
rect 21998 421 22183 427
rect 21616 370 21885 384
rect -237 359 -171 365
rect 2391 361 2457 370
rect 5629 361 5695 370
rect 8867 361 8933 370
rect 12105 361 12171 370
rect 15343 361 15409 370
rect 18581 361 18647 370
rect 21819 361 21885 370
rect 2391 355 2647 361
rect 2391 301 2581 355
rect 2635 301 2647 355
rect 5629 355 5885 361
rect 2391 295 2647 301
rect 5629 301 5819 355
rect 5873 301 5885 355
rect 8867 355 9123 361
rect 5629 295 5885 301
rect 8867 301 9057 355
rect 9111 301 9123 355
rect 12105 355 12361 361
rect 8867 295 9123 301
rect 12105 301 12295 355
rect 12349 301 12361 355
rect 15343 355 15599 361
rect 12105 295 12361 301
rect 15343 301 15533 355
rect 15587 301 15599 355
rect 18581 355 18837 361
rect 15343 295 15599 301
rect 18581 301 18771 355
rect 18825 301 18837 355
rect 21819 355 22075 361
rect 18581 295 18837 301
rect 21819 301 22009 355
rect 22063 301 22075 355
rect 21819 295 22075 301
rect -237 287 -171 293
<< via1 >>
rect 413 531 479 597
rect 2555 523 2621 589
rect 3651 531 3717 597
rect 5810 521 5876 587
rect 6889 531 6955 597
rect 9046 521 9112 587
rect 10127 531 10193 597
rect 12286 521 12352 587
rect 13365 531 13431 597
rect 15522 521 15588 587
rect 16603 531 16669 597
rect 18762 521 18828 587
rect 19841 531 19907 597
rect 21998 521 22064 587
rect -136 454 -84 460
rect -136 414 -130 454
rect -130 414 -90 454
rect -90 414 -84 454
rect -136 408 -84 414
rect 1010 374 1062 426
rect 4248 374 4300 426
rect 7486 374 7538 426
rect 10724 374 10776 426
rect 13962 374 14014 426
rect 17200 374 17252 426
rect 20438 374 20490 426
rect 23678 374 23730 426
rect -237 353 -171 359
rect -237 299 -231 353
rect -231 299 -177 353
rect -177 299 -171 353
rect 1738 306 1792 358
rect -237 293 -171 299
rect 4976 306 5030 358
rect 8214 306 8268 358
rect 11452 306 11506 358
rect 14690 306 14744 358
rect 17928 306 17982 358
rect 21166 306 21220 358
rect 24406 306 24460 358
<< metal2 >>
rect 412 687 2622 753
rect 3650 687 5876 753
rect 6888 687 9112 753
rect 10126 687 12352 753
rect 13364 687 15588 753
rect 16602 687 18828 753
rect 19840 687 22064 753
rect 413 597 479 687
rect 413 525 479 531
rect 2555 589 2621 687
rect 3651 597 3717 687
rect 3651 525 3717 531
rect 5810 587 5876 687
rect 2555 517 2621 523
rect 6889 597 6955 687
rect 6889 525 6955 531
rect 9046 587 9112 687
rect 5810 515 5876 521
rect 10127 597 10193 687
rect 10127 525 10193 531
rect 12286 587 12352 687
rect 9046 515 9112 521
rect 13365 597 13431 687
rect 13365 525 13431 531
rect 15522 587 15588 687
rect 12286 515 12352 521
rect 16603 597 16669 687
rect 16603 525 16669 531
rect 18762 587 18828 687
rect 15522 515 15588 521
rect 19841 597 19907 687
rect 19841 525 19907 531
rect 21998 587 22064 687
rect 18762 515 18828 521
rect 21998 515 22064 521
rect -142 408 -136 460
rect -84 458 -78 460
rect 1018 458 3340 468
rect 9722 460 9816 468
rect 16198 460 16292 468
rect 7494 458 9816 460
rect 13970 458 16292 460
rect 20446 458 22754 460
rect -84 410 434 458
rect 1018 432 3672 458
rect 6484 448 6910 458
rect 4252 432 6910 448
rect 7494 432 10148 458
rect 12960 448 13386 458
rect 10728 432 13386 448
rect 13970 432 16624 458
rect 19436 448 19862 458
rect 17204 432 19862 448
rect 20446 432 23102 458
rect -84 408 -78 410
rect 386 374 434 410
rect 1004 426 3672 432
rect 1004 374 1010 426
rect 1062 420 3672 426
rect 1062 374 1070 420
rect 3246 410 3672 420
rect -236 359 -172 362
rect -243 293 -237 359
rect -171 293 5 359
rect 386 326 1070 374
rect 3624 374 3672 410
rect 4242 426 6910 432
rect 4242 374 4248 426
rect 4300 410 6910 426
rect 4300 400 6568 410
rect 4300 374 4308 400
rect 1730 358 1796 366
rect -236 288 -172 293
rect -61 261 5 293
rect 1730 306 1738 358
rect 1792 306 1796 358
rect 3624 326 4308 374
rect 6862 374 6910 410
rect 7480 426 10148 432
rect 7480 374 7486 426
rect 7538 412 10148 426
rect 7538 374 7546 412
rect 9722 410 10148 412
rect 4968 358 5034 366
rect 1730 261 1796 306
rect 4968 306 4976 358
rect 5030 306 5034 358
rect 6862 326 7546 374
rect 10100 374 10148 410
rect 10718 426 13386 432
rect 10718 374 10724 426
rect 10776 410 13386 426
rect 10776 400 13044 410
rect 10776 374 10784 400
rect 8206 358 8272 366
rect 4968 261 5034 306
rect 8206 306 8214 358
rect 8268 306 8272 358
rect 10100 326 10784 374
rect 13338 374 13386 410
rect 13956 426 16624 432
rect 13956 374 13962 426
rect 14014 412 16624 426
rect 14014 374 14022 412
rect 16198 410 16624 412
rect 11444 358 11510 366
rect 8206 261 8272 306
rect 11444 306 11452 358
rect 11506 306 11510 358
rect 13338 326 14022 374
rect 16576 374 16624 410
rect 17194 426 19862 432
rect 17194 374 17200 426
rect 17252 410 19862 426
rect 17252 400 19520 410
rect 17252 374 17260 400
rect 14682 358 14748 366
rect 11444 261 11510 306
rect 14682 306 14690 358
rect 14744 306 14748 358
rect 16576 326 17260 374
rect 19814 374 19862 410
rect 20432 426 23102 432
rect 20432 374 20438 426
rect 20490 412 23102 426
rect 20490 374 20498 412
rect 22656 410 23102 412
rect 17920 358 17986 366
rect 14682 261 14748 306
rect 17920 306 17928 358
rect 17982 306 17986 358
rect 19814 326 20498 374
rect 23054 374 23102 410
rect 23672 426 23738 432
rect 23672 374 23678 426
rect 23730 374 23738 426
rect 21158 358 21224 366
rect 17920 261 17986 306
rect 21158 306 21166 358
rect 21220 306 21224 358
rect 23054 326 23738 374
rect 24398 358 24464 366
rect 21158 261 21224 306
rect 24398 306 24406 358
rect 24460 306 24464 358
rect 22650 261 22692 262
rect 24398 261 24464 306
rect -61 195 24464 261
rect 22650 194 22692 195
use inv  inv_0 ~/magic/library/mag
timestamp 1738780557
transform 1 0 22352 0 1 0
box -4 0 322 976
use inv  inv_1
timestamp 1738780557
transform 1 0 -314 0 1 0
box -4 0 322 976
use inv  inv_2
timestamp 1738780557
transform 1 0 2924 0 1 0
box -4 0 322 976
use inv  inv_3
timestamp 1738780557
transform 1 0 6162 0 1 0
box -4 0 322 976
use inv  inv_4
timestamp 1738780557
transform 1 0 9400 0 1 0
box -4 0 322 976
use inv  inv_5
timestamp 1738780557
transform 1 0 19114 0 1 0
box -4 0 322 976
use inv  inv_6
timestamp 1738780557
transform 1 0 15876 0 1 0
box -4 0 322 976
use inv  inv_7
timestamp 1738780557
transform 1 0 12638 0 1 0
box -4 0 322 976
use nand  nand_0 ~/magic/library/mag
timestamp 1739944168
transform 1 0 8974 0 1 0
box -4 0 430 976
use nand  nand_1
timestamp 1739944168
transform 1 0 2498 0 1 0
box -4 0 430 976
use nand  nand_2
timestamp 1739944168
transform 1 0 5736 0 1 0
box -4 0 430 976
use nand  nand_3
timestamp 1739944168
transform 1 0 21926 0 1 0
box -4 0 430 976
use nand  nand_4
timestamp 1739944168
transform 1 0 18688 0 1 0
box -4 0 430 976
use nand  nand_5
timestamp 1739944168
transform 1 0 15450 0 1 0
box -4 0 430 976
use nand  nand_6
timestamp 1739944168
transform 1 0 12212 0 1 0
box -4 0 430 976
use tff  tff_0
timestamp 1745480928
transform 1 0 6776 0 1 0
box -300 0 2212 976
use tff  tff_1
timestamp 1745480928
transform 1 0 300 0 1 0
box -300 0 2212 976
use tff  tff_2
timestamp 1745480928
transform 1 0 3538 0 1 0
box -300 0 2212 976
use tff  tff_3
timestamp 1745480928
transform 1 0 22968 0 1 0
box -300 0 2212 976
use tff  tff_4
timestamp 1745480928
transform 1 0 10014 0 1 0
box -300 0 2212 976
use tff  tff_5
timestamp 1745480928
transform 1 0 19728 0 1 0
box -300 0 2212 976
use tff  tff_6
timestamp 1745480928
transform 1 0 16490 0 1 0
box -300 0 2212 976
use tff  tff_7
timestamp 1745480928
transform 1 0 13252 0 1 0
box -300 0 2212 976
<< labels >>
flabel metal2 -236 288 -172 362 0 FreeSerif 160 0 0 0 CLK
port 2 nsew
flabel metal1 2391 296 2502 360 0 FreeSerif 160 0 0 0 Q0
port 5 nsew
flabel metal1 5630 296 5774 360 0 FreeSerif 160 0 0 0 Q1
port 9 nsew
flabel metal1 8870 296 9008 360 0 FreeSerif 160 0 0 0 Q2
port 13 nsew
flabel locali -314 864 22674 960 0 FreeSerif 160 0 0 0 VDD!
flabel locali -314 0 22674 96 0 FreeSerif 160 0 0 0 GND!
flabel metal1 12106 296 12250 360 0 FreeSerif 160 0 0 0 Q3
port 17 nsew
flabel metal1 15346 296 15484 360 0 FreeSerif 160 0 0 0 Q4
port 21 nsew
flabel metal1 18582 296 18726 360 0 FreeSerif 160 0 0 0 Q5
port 25 nsew
flabel metal1 21822 296 21960 360 0 FreeSerif 160 0 0 0 Q6
port 29 nsew
flabel locali 24856 370 24922 436 0 FreeSerif 160 0 0 0 Q7
port 32 nsew
<< end >>
