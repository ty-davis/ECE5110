magic
tech sky130A
timestamp 1744679307
<< poly >>
rect -51 -17 996 0
rect -51 -88 996 -71
rect -51 -159 996 -142
rect -51 -230 996 -213
rect -51 -301 996 -284
rect -51 -372 996 -355
rect -51 -443 996 -426
rect -51 -514 996 -497
rect -51 -585 996 -568
rect -51 -656 996 -639
rect -51 -727 996 -710
rect -51 -798 996 -781
rect -51 -869 996 -852
rect -51 -940 996 -923
rect -51 -1011 996 -994
rect -51 -1082 996 -1065
rect -51 -1153 996 -1136
rect -51 -1224 996 -1207
rect -51 -1295 996 -1278
rect -51 -1366 996 -1349
rect -51 -1437 996 -1420
rect -51 -1508 996 -1491
rect -51 -1579 996 -1562
rect -51 -1650 996 -1633
rect -51 -1721 996 -1704
rect -51 -1792 996 -1775
rect -51 -1863 996 -1846
rect -51 -1934 996 -1917
rect -51 -2005 996 -1988
rect -51 -2076 996 -2059
rect -51 -2147 996 -2130
rect -51 -2218 996 -2201
rect -51 -2289 996 -2272
rect -51 -2360 996 -2343
rect -51 -2431 996 -2414
rect -51 -2502 996 -2485
rect -51 -2573 996 -2556
rect -51 -2644 996 -2627
rect -51 -2715 996 -2698
rect -51 -2786 996 -2769
rect -51 -2857 996 -2840
rect -51 -2928 996 -2911
rect -51 -2999 996 -2982
rect -51 -3070 996 -3053
rect -51 -3141 996 -3124
rect -51 -3212 996 -3195
rect -51 -3283 996 -3266
rect -51 -3354 996 -3337
rect -51 -3425 996 -3408
rect -51 -3496 996 -3479
rect -51 -3567 996 -3550
rect -51 -3638 996 -3621
rect -51 -3709 996 -3692
rect -51 -3780 996 -3763
rect -51 -3851 996 -3834
rect -51 -3922 996 -3905
rect -51 -3993 996 -3976
rect -51 -4064 996 -4047
rect -51 -4135 996 -4118
rect -51 -4206 996 -4189
rect -51 -4277 996 -4260
rect -51 -4348 996 -4331
rect -51 -4419 996 -4402
rect -51 -4490 996 -4473
rect -51 -4561 996 -4544
rect -51 -4632 996 -4615
rect -51 -4703 996 -4686
rect -51 -4774 996 -4757
rect -51 -4845 996 -4828
rect -51 -4916 996 -4899
rect -51 -4987 996 -4970
rect -51 -5058 996 -5041
rect -51 -5129 996 -5112
rect -51 -5200 996 -5183
rect -51 -5271 996 -5254
rect -51 -5342 996 -5325
rect -51 -5413 996 -5396
rect -51 -5484 996 -5467
rect -51 -5555 996 -5538
rect -51 -5626 996 -5609
rect -51 -5697 996 -5680
rect -51 -5768 996 -5751
rect -51 -5839 996 -5822
rect -51 -5910 996 -5893
rect -51 -5981 996 -5964
rect -51 -6052 996 -6035
rect -51 -6123 996 -6106
rect -51 -6194 996 -6177
rect -51 -6265 996 -6248
rect -51 -6336 996 -6319
rect -51 -6407 996 -6390
rect -51 -6478 996 -6461
rect -51 -6549 996 -6532
rect -51 -6620 996 -6603
rect -51 -6691 996 -6674
rect -51 -6762 996 -6745
rect -51 -6833 996 -6816
rect -51 -6904 996 -6887
rect -51 -6975 996 -6958
rect -51 -7046 996 -7029
rect -51 -7117 996 -7100
rect -51 -7188 996 -7171
rect -51 -7259 996 -7242
rect -51 -7330 996 -7313
rect -51 -7401 996 -7384
rect -51 -7472 996 -7455
rect -51 -7543 996 -7526
rect -51 -7614 996 -7597
rect -51 -7685 996 -7668
rect -51 -7756 996 -7739
rect -51 -7827 996 -7810
rect -51 -7898 996 -7881
rect -51 -7969 996 -7952
rect -51 -8040 996 -8023
rect -51 -8111 996 -8094
rect -51 -8182 996 -8165
rect -51 -8253 996 -8236
rect -51 -8324 996 -8307
rect -51 -8395 996 -8378
rect -51 -8466 996 -8449
rect -51 -8537 996 -8520
rect -51 -8608 996 -8591
rect -51 -8679 996 -8662
rect -51 -8750 996 -8733
rect -51 -8821 996 -8804
rect -51 -8892 996 -8875
rect -51 -8963 996 -8946
rect -51 -9034 996 -9017
<< locali >>
rect 0 -9088 33 41
rect 83 -9088 116 41
rect 166 -9088 199 41
rect 249 -9088 282 41
rect 332 -9088 365 41
rect 415 -9088 448 41
rect 498 -9088 531 41
rect 581 -9088 614 41
rect 664 -9088 697 41
rect 747 -9088 780 41
rect 830 -9088 863 41
rect 913 -9088 946 41
<< ndiff >>
rect 116 -1196 208 -1163
rect 614 -1196 706 -1163
rect -9 -1196 83 -1163
rect 83 -1196 116 -1163
rect 830 -1196 863 -1163
rect 240 -1196 332 -1163
rect 581 -1196 614 -1163
rect 738 -1196 830 -1163
rect 365 -1196 457 -1163
rect 489 -1196 581 -1163
rect 332 -1196 365 -1163
rect 863 -1196 955 -1163
rect 116 -1338 208 -1305
rect 614 -1338 706 -1305
rect -9 -1338 83 -1305
rect 83 -1338 116 -1305
rect 830 -1338 863 -1305
rect 240 -1338 332 -1305
rect 581 -1338 614 -1305
rect 738 -1338 830 -1305
rect 365 -1338 457 -1305
rect 489 -1338 581 -1305
rect 332 -1338 365 -1305
rect 863 -1338 955 -1305
rect 116 -1480 208 -1447
rect 614 -1480 706 -1447
rect -9 -1480 83 -1447
rect 83 -1480 116 -1447
rect 830 -1480 863 -1447
rect 240 -1480 332 -1447
rect 581 -1480 614 -1447
rect 738 -1480 830 -1447
rect 365 -1480 457 -1447
rect 489 -1480 581 -1447
rect 332 -1480 365 -1447
rect 863 -1480 955 -1447
rect 116 -1622 208 -1589
rect 614 -1622 706 -1589
rect -9 -1622 83 -1589
rect 83 -1622 116 -1589
rect 830 -1622 863 -1589
rect 240 -1622 332 -1589
rect 581 -1622 614 -1589
rect 738 -1622 830 -1589
rect 365 -1622 457 -1589
rect 489 -1622 581 -1589
rect 332 -1622 365 -1589
rect 863 -1622 955 -1589
rect 116 -1764 208 -1731
rect 614 -1764 706 -1731
rect -9 -1764 83 -1731
rect 83 -1764 116 -1731
rect 830 -1764 863 -1731
rect 240 -1764 332 -1731
rect 581 -1764 614 -1731
rect 738 -1764 830 -1731
rect 365 -1764 457 -1731
rect 489 -1764 581 -1731
rect 332 -1764 365 -1731
rect 863 -1764 955 -1731
rect 116 -1906 208 -1873
rect 614 -1906 706 -1873
rect -9 -1906 83 -1873
rect 83 -1906 116 -1873
rect 830 -1906 863 -1873
rect 240 -1906 332 -1873
rect 581 -1906 614 -1873
rect 738 -1906 830 -1873
rect 365 -1906 457 -1873
rect 489 -1906 581 -1873
rect 332 -1906 365 -1873
rect 863 -1906 955 -1873
rect 116 -2048 208 -2015
rect 614 -2048 706 -2015
rect -9 -2048 83 -2015
rect 83 -2048 116 -2015
rect 830 -2048 863 -2015
rect 240 -2048 332 -2015
rect 581 -2048 614 -2015
rect 738 -2048 830 -2015
rect 365 -2048 457 -2015
rect 489 -2048 581 -2015
rect 332 -2048 365 -2015
rect 863 -2048 955 -2015
rect 116 -2190 208 -2157
rect 614 -2190 706 -2157
rect -9 -2190 83 -2157
rect 83 -2190 116 -2157
rect 830 -2190 863 -2157
rect 240 -2190 332 -2157
rect 581 -2190 614 -2157
rect 738 -2190 830 -2157
rect 365 -2190 457 -2157
rect 489 -2190 581 -2157
rect 332 -2190 365 -2157
rect 863 -2190 955 -2157
rect 614 -2332 706 -2299
rect 830 -2332 863 -2299
rect 581 -2332 614 -2299
rect 738 -2332 830 -2299
rect 489 -2332 581 -2299
rect 863 -2332 955 -2299
rect 614 -2474 706 -2441
rect 830 -2474 863 -2441
rect 240 -2474 332 -2441
rect 581 -2474 614 -2441
rect 738 -2474 830 -2441
rect 365 -2474 457 -2441
rect 489 -2474 581 -2441
rect 332 -2474 365 -2441
rect 863 -2474 955 -2441
rect 116 -2616 208 -2583
rect 614 -2616 706 -2583
rect 83 -2616 116 -2583
rect 830 -2616 863 -2583
rect 240 -2616 332 -2583
rect 581 -2616 614 -2583
rect 738 -2616 830 -2583
rect 365 -2616 457 -2583
rect 489 -2616 581 -2583
rect 332 -2616 365 -2583
rect 863 -2616 955 -2583
rect 116 -2758 208 -2725
rect 614 -2758 706 -2725
rect 83 -2758 116 -2725
rect 830 -2758 863 -2725
rect 240 -2758 332 -2725
rect 581 -2758 614 -2725
rect 738 -2758 830 -2725
rect 365 -2758 457 -2725
rect 489 -2758 581 -2725
rect 332 -2758 365 -2725
rect 863 -2758 955 -2725
rect 116 -2900 208 -2867
rect 614 -2900 706 -2867
rect -9 -2900 83 -2867
rect 83 -2900 116 -2867
rect 830 -2900 863 -2867
rect 240 -2900 332 -2867
rect 581 -2900 614 -2867
rect 738 -2900 830 -2867
rect 365 -2900 457 -2867
rect 489 -2900 581 -2867
rect 332 -2900 365 -2867
rect 863 -2900 955 -2867
rect 614 -3042 706 -3009
rect -9 -3042 83 -3009
rect 83 -3042 116 -3009
rect 830 -3042 863 -3009
rect 240 -3042 332 -3009
rect 581 -3042 614 -3009
rect 738 -3042 830 -3009
rect 365 -3042 457 -3009
rect 489 -3042 581 -3009
rect 332 -3042 365 -3009
rect 863 -3042 955 -3009
rect 116 -3184 208 -3151
rect 614 -3184 706 -3151
rect -9 -3184 83 -3151
rect 83 -3184 116 -3151
rect 830 -3184 863 -3151
rect 240 -3184 332 -3151
rect 581 -3184 614 -3151
rect 738 -3184 830 -3151
rect 365 -3184 457 -3151
rect 489 -3184 581 -3151
rect 332 -3184 365 -3151
rect 863 -3184 955 -3151
rect 116 -3326 208 -3293
rect 614 -3326 706 -3293
rect -9 -3326 83 -3293
rect 83 -3326 116 -3293
rect 830 -3326 863 -3293
rect 240 -3326 332 -3293
rect 581 -3326 614 -3293
rect 738 -3326 830 -3293
rect 365 -3326 457 -3293
rect 489 -3326 581 -3293
rect 332 -3326 365 -3293
rect 863 -3326 955 -3293
rect 116 -3468 208 -3435
rect 614 -3468 706 -3435
rect -9 -3468 83 -3435
rect 83 -3468 116 -3435
rect 830 -3468 863 -3435
rect 240 -3468 332 -3435
rect 581 -3468 614 -3435
rect 738 -3468 830 -3435
rect 365 -3468 457 -3435
rect 489 -3468 581 -3435
rect 332 -3468 365 -3435
rect 863 -3468 955 -3435
rect 116 -3610 208 -3577
rect 614 -3610 706 -3577
rect -9 -3610 83 -3577
rect 83 -3610 116 -3577
rect 830 -3610 863 -3577
rect 581 -3610 614 -3577
rect 738 -3610 830 -3577
rect 365 -3610 457 -3577
rect 489 -3610 581 -3577
rect 332 -3610 365 -3577
rect 863 -3610 955 -3577
rect 614 -3752 706 -3719
rect -9 -3752 83 -3719
rect 83 -3752 116 -3719
rect 830 -3752 863 -3719
rect 240 -3752 332 -3719
rect 581 -3752 614 -3719
rect 738 -3752 830 -3719
rect 365 -3752 457 -3719
rect 489 -3752 581 -3719
rect 332 -3752 365 -3719
rect 863 -3752 955 -3719
rect 614 -3894 706 -3861
rect -9 -3894 83 -3861
rect 83 -3894 116 -3861
rect 830 -3894 863 -3861
rect 581 -3894 614 -3861
rect 738 -3894 830 -3861
rect 365 -3894 457 -3861
rect 489 -3894 581 -3861
rect 332 -3894 365 -3861
rect 863 -3894 955 -3861
rect 116 -4036 208 -4003
rect 614 -4036 706 -4003
rect 83 -4036 116 -4003
rect 830 -4036 863 -4003
rect 240 -4036 332 -4003
rect 581 -4036 614 -4003
rect 738 -4036 830 -4003
rect 365 -4036 457 -4003
rect 489 -4036 581 -4003
rect 332 -4036 365 -4003
rect 863 -4036 955 -4003
rect 116 -4178 208 -4145
rect 614 -4178 706 -4145
rect 83 -4178 116 -4145
rect 830 -4178 863 -4145
rect 581 -4178 614 -4145
rect 738 -4178 830 -4145
rect 365 -4178 457 -4145
rect 489 -4178 581 -4145
rect 332 -4178 365 -4145
rect 863 -4178 955 -4145
rect 614 -4320 706 -4287
rect 830 -4320 863 -4287
rect 240 -4320 332 -4287
rect 581 -4320 614 -4287
rect 738 -4320 830 -4287
rect 365 -4320 457 -4287
rect 489 -4320 581 -4287
rect 332 -4320 365 -4287
rect 863 -4320 955 -4287
rect 614 -4462 706 -4429
rect 830 -4462 863 -4429
rect 581 -4462 614 -4429
rect 738 -4462 830 -4429
rect 365 -4462 457 -4429
rect 489 -4462 581 -4429
rect 332 -4462 365 -4429
rect 863 -4462 955 -4429
rect 614 -4604 706 -4571
rect 830 -4604 863 -4571
rect 581 -4604 614 -4571
rect 738 -4604 830 -4571
rect 863 -4604 955 -4571
rect 614 -4746 706 -4713
rect 830 -4746 863 -4713
rect 581 -4746 614 -4713
rect 738 -4746 830 -4713
rect 365 -4746 457 -4713
rect 489 -4746 581 -4713
rect 332 -4746 365 -4713
rect 863 -4746 955 -4713
rect 614 -4888 706 -4855
rect 830 -4888 863 -4855
rect 240 -4888 332 -4855
rect 581 -4888 614 -4855
rect 738 -4888 830 -4855
rect 365 -4888 457 -4855
rect 489 -4888 581 -4855
rect 332 -4888 365 -4855
rect 863 -4888 955 -4855
rect 614 -5030 706 -4997
rect 830 -5030 863 -4997
rect 240 -5030 332 -4997
rect 581 -5030 614 -4997
rect 738 -5030 830 -4997
rect 365 -5030 457 -4997
rect 489 -5030 581 -4997
rect 332 -5030 365 -4997
rect 863 -5030 955 -4997
rect 116 -5172 208 -5139
rect 614 -5172 706 -5139
rect 83 -5172 116 -5139
rect 830 -5172 863 -5139
rect 240 -5172 332 -5139
rect 581 -5172 614 -5139
rect 738 -5172 830 -5139
rect 365 -5172 457 -5139
rect 489 -5172 581 -5139
rect 332 -5172 365 -5139
rect 863 -5172 955 -5139
rect 116 -5314 208 -5281
rect 614 -5314 706 -5281
rect 83 -5314 116 -5281
rect 830 -5314 863 -5281
rect 581 -5314 614 -5281
rect 738 -5314 830 -5281
rect 365 -5314 457 -5281
rect 489 -5314 581 -5281
rect 332 -5314 365 -5281
rect 863 -5314 955 -5281
rect 116 -5456 208 -5423
rect 614 -5456 706 -5423
rect 83 -5456 116 -5423
rect 830 -5456 863 -5423
rect 240 -5456 332 -5423
rect 581 -5456 614 -5423
rect 738 -5456 830 -5423
rect 365 -5456 457 -5423
rect 489 -5456 581 -5423
rect 332 -5456 365 -5423
rect 863 -5456 955 -5423
rect 116 -5598 208 -5565
rect 614 -5598 706 -5565
rect 83 -5598 116 -5565
rect 830 -5598 863 -5565
rect 240 -5598 332 -5565
rect 581 -5598 614 -5565
rect 738 -5598 830 -5565
rect 365 -5598 457 -5565
rect 489 -5598 581 -5565
rect 332 -5598 365 -5565
rect 863 -5598 955 -5565
rect 116 -5740 208 -5707
rect 614 -5740 706 -5707
rect -9 -5740 83 -5707
rect 83 -5740 116 -5707
rect 830 -5740 863 -5707
rect 240 -5740 332 -5707
rect 581 -5740 614 -5707
rect 738 -5740 830 -5707
rect 365 -5740 457 -5707
rect 489 -5740 581 -5707
rect 332 -5740 365 -5707
rect 863 -5740 955 -5707
rect 614 -5882 706 -5849
rect -9 -5882 83 -5849
rect 83 -5882 116 -5849
rect 830 -5882 863 -5849
rect 581 -5882 614 -5849
rect 738 -5882 830 -5849
rect 365 -5882 457 -5849
rect 489 -5882 581 -5849
rect 332 -5882 365 -5849
rect 863 -5882 955 -5849
rect 614 -6024 706 -5991
rect -9 -6024 83 -5991
rect 83 -6024 116 -5991
rect 830 -6024 863 -5991
rect 240 -6024 332 -5991
rect 581 -6024 614 -5991
rect 738 -6024 830 -5991
rect 365 -6024 457 -5991
rect 489 -6024 581 -5991
rect 332 -6024 365 -5991
rect 863 -6024 955 -5991
rect 614 -6166 706 -6133
rect -9 -6166 83 -6133
rect 83 -6166 116 -6133
rect 830 -6166 863 -6133
rect 240 -6166 332 -6133
rect 581 -6166 614 -6133
rect 738 -6166 830 -6133
rect 365 -6166 457 -6133
rect 489 -6166 581 -6133
rect 332 -6166 365 -6133
rect 863 -6166 955 -6133
rect 116 -6308 208 -6275
rect 614 -6308 706 -6275
rect -9 -6308 83 -6275
rect 83 -6308 116 -6275
rect 830 -6308 863 -6275
rect 240 -6308 332 -6275
rect 581 -6308 614 -6275
rect 738 -6308 830 -6275
rect 365 -6308 457 -6275
rect 489 -6308 581 -6275
rect 332 -6308 365 -6275
rect 863 -6308 955 -6275
rect 116 -6450 208 -6417
rect 614 -6450 706 -6417
rect -9 -6450 83 -6417
rect 83 -6450 116 -6417
rect 830 -6450 863 -6417
rect 581 -6450 614 -6417
rect 738 -6450 830 -6417
rect 365 -6450 457 -6417
rect 489 -6450 581 -6417
rect 332 -6450 365 -6417
rect 863 -6450 955 -6417
rect 116 -6592 208 -6559
rect 614 -6592 706 -6559
rect -9 -6592 83 -6559
rect 83 -6592 116 -6559
rect 830 -6592 863 -6559
rect 240 -6592 332 -6559
rect 581 -6592 614 -6559
rect 738 -6592 830 -6559
rect 365 -6592 457 -6559
rect 489 -6592 581 -6559
rect 332 -6592 365 -6559
rect 863 -6592 955 -6559
rect 116 -6734 208 -6701
rect 614 -6734 706 -6701
rect -9 -6734 83 -6701
rect 83 -6734 116 -6701
rect 830 -6734 863 -6701
rect 240 -6734 332 -6701
rect 581 -6734 614 -6701
rect 738 -6734 830 -6701
rect 365 -6734 457 -6701
rect 489 -6734 581 -6701
rect 332 -6734 365 -6701
rect 863 -6734 955 -6701
rect 830 -6876 863 -6843
rect 738 -6876 830 -6843
rect 614 -7018 706 -6985
rect 830 -7018 863 -6985
rect 581 -7018 614 -6985
rect 738 -7018 830 -6985
rect 365 -7018 457 -6985
rect 489 -7018 581 -6985
rect 332 -7018 365 -6985
rect 863 -7018 955 -6985
rect 614 -7160 706 -7127
rect 830 -7160 863 -7127
rect 240 -7160 332 -7127
rect 581 -7160 614 -7127
rect 365 -7160 457 -7127
rect 489 -7160 581 -7127
rect 332 -7160 365 -7127
rect 863 -7160 955 -7127
rect 116 -7302 208 -7269
rect 614 -7302 706 -7269
rect 83 -7302 116 -7269
rect 830 -7302 863 -7269
rect 240 -7302 332 -7269
rect 581 -7302 614 -7269
rect 738 -7302 830 -7269
rect 489 -7302 581 -7269
rect 332 -7302 365 -7269
rect 863 -7302 955 -7269
rect -9 -7444 83 -7411
rect 83 -7444 116 -7411
rect 581 -7444 614 -7411
rect 365 -7444 457 -7411
rect 489 -7444 581 -7411
rect 332 -7444 365 -7411
rect 116 -7586 208 -7553
rect -9 -7586 83 -7553
rect 614 -7586 706 -7553
rect 83 -7586 116 -7553
rect 830 -7586 863 -7553
rect 240 -7586 332 -7553
rect 581 -7586 614 -7553
rect 365 -7586 457 -7553
rect 738 -7586 830 -7553
rect 332 -7586 365 -7553
rect 116 -7728 208 -7695
rect -9 -7728 83 -7695
rect 83 -7728 116 -7695
rect 830 -7728 863 -7695
rect 240 -7728 332 -7695
rect 581 -7728 614 -7695
rect 738 -7728 830 -7695
rect 365 -7728 457 -7695
rect 489 -7728 581 -7695
rect 332 -7728 365 -7695
rect 116 -7870 208 -7837
rect 614 -7870 706 -7837
rect -9 -7870 83 -7837
rect 83 -7870 116 -7837
rect 830 -7870 863 -7837
rect 240 -7870 332 -7837
rect 581 -7870 614 -7837
rect 365 -7870 457 -7837
rect 489 -7870 581 -7837
rect 332 -7870 365 -7837
rect 863 -7870 955 -7837
rect 116 -8012 208 -7979
rect 614 -8012 706 -7979
rect -9 -8012 83 -7979
rect 83 -8012 116 -7979
rect 830 -8012 863 -7979
rect 240 -8012 332 -7979
rect 581 -8012 614 -7979
rect 738 -8012 830 -7979
rect 365 -8012 457 -7979
rect 489 -8012 581 -7979
rect 332 -8012 365 -7979
rect 863 -8012 955 -7979
rect 116 -8154 208 -8121
rect 614 -8154 706 -8121
rect -9 -8154 83 -8121
rect 83 -8154 116 -8121
rect 830 -8154 863 -8121
rect 240 -8154 332 -8121
rect 581 -8154 614 -8121
rect 365 -8154 457 -8121
rect 738 -8154 830 -8121
rect 489 -8154 581 -8121
rect 332 -8154 365 -8121
rect 863 -8154 955 -8121
rect 116 -8296 208 -8263
rect -9 -8296 83 -8263
rect 614 -8296 706 -8263
rect 83 -8296 116 -8263
rect 830 -8296 863 -8263
rect 581 -8296 614 -8263
rect 738 -8296 830 -8263
rect 365 -8296 457 -8263
rect 489 -8296 581 -8263
rect 332 -8296 365 -8263
rect -9 -8438 83 -8405
rect 83 -8438 116 -8405
rect 240 -8438 332 -8405
rect 581 -8438 614 -8405
rect 365 -8438 457 -8405
rect 489 -8438 581 -8405
rect 332 -8438 365 -8405
rect 116 -8580 208 -8547
rect -9 -8580 83 -8547
rect 614 -8580 706 -8547
rect 83 -8580 116 -8547
rect 830 -8580 863 -8547
rect 240 -8580 332 -8547
rect 581 -8580 614 -8547
rect 738 -8580 830 -8547
rect 332 -8580 365 -8547
rect 863 -8580 955 -8547
rect 116 -8722 208 -8689
rect 614 -8722 706 -8689
rect 83 -8722 116 -8689
rect 830 -8722 863 -8689
rect 240 -8722 332 -8689
rect 581 -8722 614 -8689
rect 738 -8722 830 -8689
rect 365 -8722 457 -8689
rect 489 -8722 581 -8689
rect 332 -8722 365 -8689
rect 863 -8722 955 -8689
rect 614 -8864 706 -8831
rect 830 -8864 863 -8831
rect 240 -8864 332 -8831
rect 581 -8864 614 -8831
rect 365 -8864 457 -8831
rect 332 -8864 365 -8831
rect 863 -8864 955 -8831
rect 830 -9006 863 -8973
rect 738 -9006 830 -8973
rect 489 -9006 581 -8973
rect 581 -9006 614 -8973
rect 655 -1125 706 -1092
rect 904 -1125 955 -1092
rect 489 -1125 540 -1092
rect 738 -1125 789 -1092
rect 157 -1125 208 -1092
rect 406 -1125 457 -1092
rect -9 -1125 42 -1092
rect 240 -1125 291 -1092
rect 655 -1267 706 -1234
rect 904 -1267 955 -1234
rect 489 -1267 540 -1234
rect 738 -1267 789 -1234
rect 157 -1267 208 -1234
rect 406 -1267 457 -1234
rect -9 -1267 42 -1234
rect 240 -1267 291 -1234
rect 655 -1409 706 -1376
rect 904 -1409 955 -1376
rect 489 -1409 540 -1376
rect 738 -1409 789 -1376
rect 157 -1409 208 -1376
rect 406 -1409 457 -1376
rect -9 -1409 42 -1376
rect 240 -1409 291 -1376
rect 655 -1551 706 -1518
rect 904 -1551 955 -1518
rect 489 -1551 540 -1518
rect 738 -1551 789 -1518
rect 157 -1551 208 -1518
rect 406 -1551 457 -1518
rect -9 -1551 42 -1518
rect 240 -1551 291 -1518
rect 655 -1693 706 -1660
rect 904 -1693 955 -1660
rect 489 -1693 540 -1660
rect 738 -1693 789 -1660
rect 157 -1693 208 -1660
rect 406 -1693 457 -1660
rect -9 -1693 42 -1660
rect 240 -1693 291 -1660
rect 655 -1835 706 -1802
rect 904 -1835 955 -1802
rect 489 -1835 540 -1802
rect 738 -1835 789 -1802
rect 157 -1835 208 -1802
rect 406 -1835 457 -1802
rect -9 -1835 42 -1802
rect 240 -1835 291 -1802
rect 655 -1977 706 -1944
rect 904 -1977 955 -1944
rect 489 -1977 540 -1944
rect 738 -1977 789 -1944
rect 157 -1977 208 -1944
rect 406 -1977 457 -1944
rect -9 -1977 42 -1944
rect 240 -1977 291 -1944
rect 655 -2119 706 -2086
rect 904 -2119 955 -2086
rect 489 -2119 540 -2086
rect 738 -2119 789 -2086
rect 157 -2119 208 -2086
rect 406 -2119 457 -2086
rect -9 -2119 42 -2086
rect 240 -2119 291 -2086
rect 655 -2261 706 -2228
rect 904 -2261 955 -2228
rect 489 -2261 540 -2228
rect 738 -2261 789 -2228
rect 157 -2261 208 -2228
rect 406 -2261 457 -2228
rect -9 -2261 42 -2228
rect 240 -2261 291 -2228
rect 655 -2403 706 -2370
rect 904 -2403 955 -2370
rect 489 -2403 540 -2370
rect 738 -2403 789 -2370
rect 406 -2403 457 -2370
rect 655 -2545 706 -2512
rect 904 -2545 955 -2512
rect 489 -2545 540 -2512
rect 738 -2545 789 -2512
rect 406 -2545 457 -2512
rect 240 -2545 291 -2512
rect 655 -2687 706 -2654
rect 904 -2687 955 -2654
rect 489 -2687 540 -2654
rect 738 -2687 789 -2654
rect 157 -2687 208 -2654
rect 406 -2687 457 -2654
rect 655 -2829 706 -2796
rect 904 -2829 955 -2796
rect 489 -2829 540 -2796
rect 738 -2829 789 -2796
rect 157 -2829 208 -2796
rect 406 -2829 457 -2796
rect 240 -2829 291 -2796
rect 655 -2971 706 -2938
rect 904 -2971 955 -2938
rect 489 -2971 540 -2938
rect 738 -2971 789 -2938
rect 406 -2971 457 -2938
rect -9 -2971 42 -2938
rect 655 -3113 706 -3080
rect 904 -3113 955 -3080
rect 489 -3113 540 -3080
rect 738 -3113 789 -3080
rect 406 -3113 457 -3080
rect -9 -3113 42 -3080
rect 240 -3113 291 -3080
rect 655 -3255 706 -3222
rect 904 -3255 955 -3222
rect 489 -3255 540 -3222
rect 738 -3255 789 -3222
rect 157 -3255 208 -3222
rect 406 -3255 457 -3222
rect -9 -3255 42 -3222
rect 655 -3397 706 -3364
rect 904 -3397 955 -3364
rect 489 -3397 540 -3364
rect 738 -3397 789 -3364
rect 157 -3397 208 -3364
rect 406 -3397 457 -3364
rect -9 -3397 42 -3364
rect 240 -3397 291 -3364
rect 655 -3539 706 -3506
rect 904 -3539 955 -3506
rect 489 -3539 540 -3506
rect 738 -3539 789 -3506
rect 157 -3539 208 -3506
rect 406 -3539 457 -3506
rect -9 -3539 42 -3506
rect 240 -3539 291 -3506
rect 655 -3681 706 -3648
rect 904 -3681 955 -3648
rect 489 -3681 540 -3648
rect 738 -3681 789 -3648
rect 157 -3681 208 -3648
rect 406 -3681 457 -3648
rect -9 -3681 42 -3648
rect 240 -3681 291 -3648
rect 655 -3823 706 -3790
rect 904 -3823 955 -3790
rect 489 -3823 540 -3790
rect 738 -3823 789 -3790
rect 406 -3823 457 -3790
rect -9 -3823 42 -3790
rect 240 -3823 291 -3790
rect 655 -3965 706 -3932
rect 904 -3965 955 -3932
rect 489 -3965 540 -3932
rect 738 -3965 789 -3932
rect 157 -3965 208 -3932
rect 406 -3965 457 -3932
rect -9 -3965 42 -3932
rect 240 -3965 291 -3932
rect 655 -4107 706 -4074
rect 904 -4107 955 -4074
rect 489 -4107 540 -4074
rect 738 -4107 789 -4074
rect 157 -4107 208 -4074
rect 406 -4107 457 -4074
rect 240 -4107 291 -4074
rect 655 -4249 706 -4216
rect 904 -4249 955 -4216
rect 489 -4249 540 -4216
rect 738 -4249 789 -4216
rect 157 -4249 208 -4216
rect 406 -4249 457 -4216
rect 240 -4249 291 -4216
rect 655 -4391 706 -4358
rect 904 -4391 955 -4358
rect 489 -4391 540 -4358
rect 738 -4391 789 -4358
rect 406 -4391 457 -4358
rect 240 -4391 291 -4358
rect 655 -4533 706 -4500
rect 904 -4533 955 -4500
rect 489 -4533 540 -4500
rect 738 -4533 789 -4500
rect 655 -4675 706 -4642
rect 904 -4675 955 -4642
rect 489 -4675 540 -4642
rect 738 -4675 789 -4642
rect 655 -4817 706 -4784
rect 904 -4817 955 -4784
rect 489 -4817 540 -4784
rect 738 -4817 789 -4784
rect 406 -4817 457 -4784
rect 655 -4959 706 -4926
rect 904 -4959 955 -4926
rect 489 -4959 540 -4926
rect 738 -4959 789 -4926
rect 240 -4959 291 -4926
rect 655 -5101 706 -5068
rect 904 -5101 955 -5068
rect 489 -5101 540 -5068
rect 738 -5101 789 -5068
rect 406 -5101 457 -5068
rect 240 -5101 291 -5068
rect 655 -5243 706 -5210
rect 904 -5243 955 -5210
rect 489 -5243 540 -5210
rect 738 -5243 789 -5210
rect 157 -5243 208 -5210
rect 655 -5385 706 -5352
rect 904 -5385 955 -5352
rect 489 -5385 540 -5352
rect 738 -5385 789 -5352
rect 157 -5385 208 -5352
rect 406 -5385 457 -5352
rect 655 -5527 706 -5494
rect 904 -5527 955 -5494
rect 489 -5527 540 -5494
rect 738 -5527 789 -5494
rect 157 -5527 208 -5494
rect 240 -5527 291 -5494
rect 655 -5669 706 -5636
rect 904 -5669 955 -5636
rect 489 -5669 540 -5636
rect 738 -5669 789 -5636
rect 157 -5669 208 -5636
rect 406 -5669 457 -5636
rect 240 -5669 291 -5636
rect 655 -5811 706 -5778
rect 904 -5811 955 -5778
rect 489 -5811 540 -5778
rect 738 -5811 789 -5778
rect -9 -5811 42 -5778
rect 655 -5953 706 -5920
rect 904 -5953 955 -5920
rect 489 -5953 540 -5920
rect 738 -5953 789 -5920
rect 406 -5953 457 -5920
rect -9 -5953 42 -5920
rect 655 -6095 706 -6062
rect 904 -6095 955 -6062
rect 489 -6095 540 -6062
rect 738 -6095 789 -6062
rect -9 -6095 42 -6062
rect 240 -6095 291 -6062
rect 655 -6237 706 -6204
rect 904 -6237 955 -6204
rect 489 -6237 540 -6204
rect 738 -6237 789 -6204
rect 406 -6237 457 -6204
rect -9 -6237 42 -6204
rect 240 -6237 291 -6204
rect 655 -6379 706 -6346
rect 904 -6379 955 -6346
rect 489 -6379 540 -6346
rect 738 -6379 789 -6346
rect 157 -6379 208 -6346
rect -9 -6379 42 -6346
rect 655 -6521 706 -6488
rect 904 -6521 955 -6488
rect 489 -6521 540 -6488
rect 738 -6521 789 -6488
rect 157 -6521 208 -6488
rect 406 -6521 457 -6488
rect -9 -6521 42 -6488
rect 655 -6663 706 -6630
rect 904 -6663 955 -6630
rect 489 -6663 540 -6630
rect 738 -6663 789 -6630
rect 157 -6663 208 -6630
rect -9 -6663 42 -6630
rect 240 -6663 291 -6630
rect 655 -6805 706 -6772
rect 904 -6805 955 -6772
rect 738 -6805 789 -6772
rect 157 -6805 208 -6772
rect 406 -6805 457 -6772
rect -9 -6805 42 -6772
rect 240 -6805 291 -6772
rect 489 -6947 540 -6914
rect 738 -6947 789 -6914
rect 655 -7089 706 -7056
rect 904 -7089 955 -7056
rect 406 -7089 457 -7056
rect 240 -7089 291 -7056
rect 655 -7231 706 -7198
rect 904 -7231 955 -7198
rect 489 -7231 540 -7198
rect 738 -7231 789 -7198
rect 157 -7231 208 -7198
rect 406 -7231 457 -7198
rect 240 -7231 291 -7198
rect 655 -7373 706 -7340
rect 904 -7373 955 -7340
rect 738 -7373 789 -7340
rect 157 -7373 208 -7340
rect -9 -7373 42 -7340
rect 240 -7373 291 -7340
rect 489 -7515 540 -7482
rect 406 -7515 457 -7482
rect -9 -7515 42 -7482
rect 240 -7515 291 -7482
rect 655 -7657 706 -7624
rect 489 -7657 540 -7624
rect 738 -7657 789 -7624
rect 157 -7657 208 -7624
rect 406 -7657 457 -7624
rect -9 -7657 42 -7624
rect 655 -7799 706 -7766
rect 904 -7799 955 -7766
rect 489 -7799 540 -7766
rect 738 -7799 789 -7766
rect 157 -7799 208 -7766
rect 406 -7799 457 -7766
rect -9 -7799 42 -7766
rect 240 -7799 291 -7766
rect 655 -7941 706 -7908
rect 904 -7941 955 -7908
rect 489 -7941 540 -7908
rect 157 -7941 208 -7908
rect 738 -7941 789 -7908
rect 406 -7941 457 -7908
rect -9 -7941 42 -7908
rect 240 -7941 291 -7908
rect 655 -8083 706 -8050
rect 904 -8083 955 -8050
rect 489 -8083 540 -8050
rect 157 -8083 208 -8050
rect 406 -8083 457 -8050
rect -9 -8083 42 -8050
rect 240 -8083 291 -8050
rect 489 -8225 540 -8192
rect 738 -8225 789 -8192
rect 157 -8225 208 -8192
rect 406 -8225 457 -8192
rect -9 -8225 42 -8192
rect 240 -8225 291 -8192
rect 655 -8367 706 -8334
rect 738 -8367 789 -8334
rect 157 -8367 208 -8334
rect 406 -8367 457 -8334
rect -9 -8367 42 -8334
rect 240 -8367 291 -8334
rect 489 -8509 540 -8476
rect 406 -8509 457 -8476
rect -9 -8509 42 -8476
rect 655 -8651 706 -8618
rect 904 -8651 955 -8618
rect 489 -8651 540 -8618
rect 738 -8651 789 -8618
rect 157 -8651 208 -8618
rect 240 -8651 291 -8618
rect 655 -8793 706 -8760
rect 904 -8793 955 -8760
rect 489 -8793 540 -8760
rect 406 -8793 457 -8760
rect 240 -8793 291 -8760
rect 655 -8935 706 -8902
rect 904 -8935 955 -8902
rect 489 -8935 540 -8902
rect 738 -8935 789 -8902
rect 406 -8935 457 -8902
rect 738 -9077 789 -9044
rect 904 -6772 955 -6734
rect 904 -2157 955 -2119
rect 904 -8831 955 -8793
rect 904 -6204 955 -6166
rect 904 -3577 955 -3539
rect 904 -2938 955 -2900
rect 904 -1944 955 -1906
rect 904 -6488 955 -6450
rect 904 -3790 955 -3752
rect 904 -5565 955 -5527
rect 904 -5494 955 -5456
rect 904 -7198 955 -7160
rect 904 -4784 955 -4746
rect 904 -5068 955 -5030
rect 904 -8121 955 -8083
rect 904 -3932 955 -3894
rect 904 -3719 955 -3681
rect 904 -4855 955 -4817
rect 904 -4713 955 -4675
rect 904 -6062 955 -6024
rect 904 -4642 955 -4604
rect 904 -1163 955 -1125
rect 904 -3293 955 -3255
rect 904 -4003 955 -3965
rect 904 -4926 955 -4888
rect 904 -6559 955 -6521
rect 904 -5920 955 -5882
rect 904 -1305 955 -1267
rect 904 -5849 955 -5811
rect 904 -8760 955 -8722
rect 904 -5210 955 -5172
rect 904 -2867 955 -2829
rect 904 -6701 955 -6663
rect 904 -6417 955 -6379
rect 904 -3861 955 -3823
rect 904 -3364 955 -3326
rect 904 -5352 955 -5314
rect 904 -1376 955 -1338
rect 904 -8618 955 -8580
rect 904 -1447 955 -1409
rect 904 -2086 955 -2048
rect 904 -4997 955 -4959
rect 904 -4145 955 -4107
rect 904 -3080 955 -3042
rect 904 -8689 955 -8651
rect 904 -4216 955 -4178
rect 904 -5636 955 -5598
rect 904 -5707 955 -5669
rect 904 -6346 955 -6308
rect 904 -6630 955 -6592
rect 904 -4074 955 -4036
rect 904 -2583 955 -2545
rect 904 -5991 955 -5953
rect 904 -8902 955 -8864
rect 904 -7269 955 -7231
rect 904 -1873 955 -1835
rect 904 -5423 955 -5385
rect 904 -2441 955 -2403
rect 904 -4500 955 -4462
rect 904 -3506 955 -3468
rect 904 -1660 955 -1622
rect 904 -8050 955 -8012
rect 904 -7837 955 -7799
rect 904 -2796 955 -2758
rect 904 -6133 955 -6095
rect 904 -1802 955 -1764
rect 904 -3435 955 -3397
rect 904 -4429 955 -4391
rect 904 -4287 955 -4249
rect 904 -3648 955 -3610
rect 904 -5139 955 -5101
rect 904 -2725 955 -2687
rect 904 -3222 955 -3184
rect 904 -7908 955 -7870
rect 904 -1234 955 -1196
rect 904 -2228 955 -2190
rect 904 -6275 955 -6237
rect 904 -5778 955 -5740
rect 904 -7979 955 -7941
rect 904 -2015 955 -1977
rect 904 -1518 955 -1480
rect 904 -3009 955 -2971
rect 904 -1589 955 -1551
rect 904 -2370 955 -2332
rect 904 -7056 955 -7018
rect 904 -7127 955 -7089
rect 904 -7340 955 -7302
rect 904 -1731 955 -1693
rect 904 -2512 955 -2474
rect 904 -3151 955 -3113
rect 904 -4358 955 -4320
rect 904 -5281 955 -5243
rect 904 -2654 955 -2616
rect 738 -6772 789 -6734
rect 738 -2157 789 -2119
rect 738 -6204 789 -6166
rect 738 -7766 789 -7728
rect 738 -3577 789 -3539
rect 738 -2938 789 -2900
rect 738 -1944 789 -1906
rect 738 -6488 789 -6450
rect 738 -3790 789 -3752
rect 738 -5565 789 -5527
rect 738 -5494 789 -5456
rect 738 -4784 789 -4746
rect 738 -5068 789 -5030
rect 738 -3932 789 -3894
rect 738 -3719 789 -3681
rect 738 -4855 789 -4817
rect 738 -4713 789 -4675
rect 738 -6062 789 -6024
rect 738 -4642 789 -4604
rect 738 -1163 789 -1125
rect 738 -3293 789 -3255
rect 738 -4003 789 -3965
rect 738 -4926 789 -4888
rect 738 -6559 789 -6521
rect 738 -5920 789 -5882
rect 738 -1305 789 -1267
rect 738 -5849 789 -5811
rect 738 -5210 789 -5172
rect 738 -2867 789 -2829
rect 738 -6701 789 -6663
rect 738 -6417 789 -6379
rect 738 -3861 789 -3823
rect 738 -3364 789 -3326
rect 738 -5352 789 -5314
rect 738 -1376 789 -1338
rect 738 -8618 789 -8580
rect 738 -1447 789 -1409
rect 738 -2086 789 -2048
rect 738 -4997 789 -4959
rect 738 -4145 789 -4107
rect 738 -3080 789 -3042
rect 738 -8689 789 -8651
rect 738 -4216 789 -4178
rect 738 -5636 789 -5598
rect 738 -7624 789 -7586
rect 738 -5707 789 -5669
rect 738 -6346 789 -6308
rect 738 -6630 789 -6592
rect 738 -4074 789 -4036
rect 738 -8263 789 -8225
rect 738 -6914 789 -6876
rect 738 -2583 789 -2545
rect 738 -5991 789 -5953
rect 738 -7269 789 -7231
rect 738 -1873 789 -1835
rect 738 -5423 789 -5385
rect 738 -9044 789 -9006
rect 738 -2441 789 -2403
rect 738 -4500 789 -4462
rect 738 -3506 789 -3468
rect 738 -1660 789 -1622
rect 738 -2796 789 -2758
rect 738 -6133 789 -6095
rect 738 -7695 789 -7657
rect 738 -1802 789 -1764
rect 738 -3435 789 -3397
rect 738 -4429 789 -4391
rect 738 -8334 789 -8296
rect 738 -4287 789 -4249
rect 738 -3648 789 -3610
rect 738 -5139 789 -5101
rect 738 -2725 789 -2687
rect 738 -3222 789 -3184
rect 738 -8973 789 -8935
rect 738 -1234 789 -1196
rect 738 -2228 789 -2190
rect 738 -6275 789 -6237
rect 738 -5778 789 -5740
rect 738 -7979 789 -7941
rect 738 -2015 789 -1977
rect 738 -1518 789 -1480
rect 738 -3009 789 -2971
rect 738 -1589 789 -1551
rect 738 -2370 789 -2332
rect 738 -7340 789 -7302
rect 738 -1731 789 -1693
rect 738 -2512 789 -2474
rect 738 -3151 789 -3113
rect 738 -4358 789 -4320
rect 738 -5281 789 -5243
rect 738 -2654 789 -2616
rect 738 -8192 789 -8154
rect 738 -6985 789 -6947
rect 655 -6772 706 -6734
rect 655 -2157 706 -2119
rect 655 -8831 706 -8793
rect 655 -6204 706 -6166
rect 655 -3577 706 -3539
rect 655 -2938 706 -2900
rect 655 -1944 706 -1906
rect 655 -6488 706 -6450
rect 655 -3790 706 -3752
rect 655 -5565 706 -5527
rect 655 -5494 706 -5456
rect 655 -4784 706 -4746
rect 655 -5068 706 -5030
rect 655 -8121 706 -8083
rect 655 -3932 706 -3894
rect 655 -3719 706 -3681
rect 655 -4855 706 -4817
rect 655 -4713 706 -4675
rect 655 -6062 706 -6024
rect 655 -4642 706 -4604
rect 655 -1163 706 -1125
rect 655 -3293 706 -3255
rect 655 -4003 706 -3965
rect 655 -4926 706 -4888
rect 655 -6559 706 -6521
rect 655 -5920 706 -5882
rect 655 -1305 706 -1267
rect 655 -5849 706 -5811
rect 655 -5210 706 -5172
rect 655 -2867 706 -2829
rect 655 -6701 706 -6663
rect 655 -6417 706 -6379
rect 655 -3861 706 -3823
rect 655 -3364 706 -3326
rect 655 -5352 706 -5314
rect 655 -1376 706 -1338
rect 655 -8618 706 -8580
rect 655 -1447 706 -1409
rect 655 -2086 706 -2048
rect 655 -4997 706 -4959
rect 655 -4145 706 -4107
rect 655 -3080 706 -3042
rect 655 -8689 706 -8651
rect 655 -4216 706 -4178
rect 655 -5636 706 -5598
rect 655 -7624 706 -7586
rect 655 -5707 706 -5669
rect 655 -6346 706 -6308
rect 655 -6630 706 -6592
rect 655 -4074 706 -4036
rect 655 -2583 706 -2545
rect 655 -5991 706 -5953
rect 655 -8902 706 -8864
rect 655 -7269 706 -7231
rect 655 -1873 706 -1835
rect 655 -5423 706 -5385
rect 655 -2441 706 -2403
rect 655 -4500 706 -4462
rect 655 -3506 706 -3468
rect 655 -1660 706 -1622
rect 655 -8050 706 -8012
rect 655 -7837 706 -7799
rect 655 -2796 706 -2758
rect 655 -6133 706 -6095
rect 655 -1802 706 -1764
rect 655 -3435 706 -3397
rect 655 -4429 706 -4391
rect 655 -8334 706 -8296
rect 655 -4287 706 -4249
rect 655 -3648 706 -3610
rect 655 -5139 706 -5101
rect 655 -2725 706 -2687
rect 655 -3222 706 -3184
rect 655 -7908 706 -7870
rect 655 -1234 706 -1196
rect 655 -2228 706 -2190
rect 655 -6275 706 -6237
rect 655 -5778 706 -5740
rect 655 -7979 706 -7941
rect 655 -2015 706 -1977
rect 655 -1518 706 -1480
rect 655 -3009 706 -2971
rect 655 -1589 706 -1551
rect 655 -2370 706 -2332
rect 655 -7056 706 -7018
rect 655 -7127 706 -7089
rect 655 -7340 706 -7302
rect 655 -1731 706 -1693
rect 655 -2512 706 -2474
rect 655 -3151 706 -3113
rect 655 -4358 706 -4320
rect 655 -5281 706 -5243
rect 655 -2654 706 -2616
rect 489 -2157 540 -2119
rect 489 -7766 540 -7728
rect 489 -3577 540 -3539
rect 489 -2938 540 -2900
rect 489 -1944 540 -1906
rect 489 -3790 540 -3752
rect 489 -5565 540 -5527
rect 489 -7198 540 -7160
rect 489 -3932 540 -3894
rect 489 -3719 540 -3681
rect 489 -4855 540 -4817
rect 489 -4713 540 -4675
rect 489 -7482 540 -7444
rect 489 -1163 540 -1125
rect 489 -3293 540 -3255
rect 489 -4003 540 -3965
rect 489 -6559 540 -6521
rect 489 -1305 540 -1267
rect 489 -5849 540 -5811
rect 489 -8476 540 -8438
rect 489 -8760 540 -8722
rect 489 -2867 540 -2829
rect 489 -6701 540 -6663
rect 489 -6417 540 -6379
rect 489 -3861 540 -3823
rect 489 -3364 540 -3326
rect 489 -1376 540 -1338
rect 489 -1447 540 -1409
rect 489 -2086 540 -2048
rect 489 -4997 540 -4959
rect 489 -4145 540 -4107
rect 489 -3080 540 -3042
rect 489 -8689 540 -8651
rect 489 -4216 540 -4178
rect 489 -5707 540 -5669
rect 489 -4074 540 -4036
rect 489 -8263 540 -8225
rect 489 -2583 540 -2545
rect 489 -5991 540 -5953
rect 489 -7269 540 -7231
rect 489 -1873 540 -1835
rect 489 -5423 540 -5385
rect 489 -2441 540 -2403
rect 489 -4500 540 -4462
rect 489 -3506 540 -3468
rect 489 -1660 540 -1622
rect 489 -8050 540 -8012
rect 489 -2796 540 -2758
rect 489 -6133 540 -6095
rect 489 -7695 540 -7657
rect 489 -1802 540 -1764
rect 489 -3435 540 -3397
rect 489 -4429 540 -4391
rect 489 -4287 540 -4249
rect 489 -3648 540 -3610
rect 489 -5139 540 -5101
rect 489 -2725 540 -2687
rect 489 -3222 540 -3184
rect 489 -8973 540 -8935
rect 489 -7908 540 -7870
rect 489 -1234 540 -1196
rect 489 -2228 540 -2190
rect 489 -6275 540 -6237
rect 489 -7979 540 -7941
rect 489 -2015 540 -1977
rect 489 -1518 540 -1480
rect 489 -3009 540 -2971
rect 489 -1589 540 -1551
rect 489 -2370 540 -2332
rect 489 -1731 540 -1693
rect 489 -2512 540 -2474
rect 489 -3151 540 -3113
rect 489 -4358 540 -4320
rect 489 -5281 540 -5243
rect 489 -2654 540 -2616
rect 489 -8192 540 -8154
rect 489 -6985 540 -6947
rect 406 -3435 457 -3397
rect 406 -4429 457 -4391
rect 406 -5920 457 -5882
rect 406 -6772 457 -6734
rect 406 -2157 457 -2119
rect 406 -4287 457 -4249
rect 406 -1305 457 -1267
rect 406 -5139 457 -5101
rect 406 -2725 457 -2687
rect 406 -6204 457 -6166
rect 406 -8476 457 -8438
rect 406 -5636 457 -5598
rect 406 -8760 457 -8722
rect 406 -7908 457 -7870
rect 406 -1234 457 -1196
rect 406 -2228 457 -2190
rect 406 -5707 457 -5669
rect 406 -3577 457 -3539
rect 406 -6275 457 -6237
rect 406 -2867 457 -2829
rect 406 -3861 457 -3823
rect 406 -8263 457 -8225
rect 406 -7979 457 -7941
rect 406 -1944 457 -1906
rect 406 -6488 457 -6450
rect 406 -7553 457 -7515
rect 406 -7198 457 -7160
rect 406 -2583 457 -2545
rect 406 -2015 457 -1977
rect 406 -4784 457 -4746
rect 406 -5068 457 -5030
rect 406 -1518 457 -1480
rect 406 -5352 457 -5314
rect 406 -5991 457 -5953
rect 406 -8121 457 -8083
rect 406 -3009 457 -2971
rect 406 -8902 457 -8864
rect 406 -3719 457 -3681
rect 406 -1873 457 -1835
rect 406 -8405 457 -8367
rect 406 -4855 457 -4817
rect 406 -5423 457 -5385
rect 406 -1376 457 -1338
rect 406 -1589 457 -1551
rect 406 -2441 457 -2403
rect 406 -1447 457 -1409
rect 406 -2086 457 -2048
rect 406 -7482 457 -7444
rect 406 -7056 457 -7018
rect 406 -1163 457 -1125
rect 406 -3293 457 -3255
rect 406 -4003 457 -3965
rect 406 -1731 457 -1693
rect 406 -4145 457 -4107
rect 406 -1660 457 -1622
rect 406 -8050 457 -8012
rect 406 -3151 457 -3113
rect 406 -7837 457 -7799
rect 406 -6559 457 -6521
rect 406 -7695 457 -7657
rect 406 -1802 457 -1764
rect 240 -3435 291 -3397
rect 240 -6772 291 -6734
rect 240 -2157 291 -2119
rect 240 -4287 291 -4249
rect 240 -1305 291 -1267
rect 240 -5139 291 -5101
rect 240 -8831 291 -8793
rect 240 -6204 291 -6166
rect 240 -7766 291 -7728
rect 240 -5636 291 -5598
rect 240 -8192 291 -8154
rect 240 -8760 291 -8722
rect 240 -7908 291 -7870
rect 240 -1234 291 -1196
rect 240 -2228 291 -2190
rect 240 -5707 291 -5669
rect 240 -6275 291 -6237
rect 240 -2867 291 -2829
rect 240 -6630 291 -6592
rect 240 -6701 291 -6663
rect 240 -4074 291 -4036
rect 240 -7979 291 -7941
rect 240 -1944 291 -1906
rect 240 -3790 291 -3752
rect 240 -7553 291 -7515
rect 240 -5565 291 -5527
rect 240 -5494 291 -5456
rect 240 -3364 291 -3326
rect 240 -7198 291 -7160
rect 240 -2583 291 -2545
rect 240 -2015 291 -1977
rect 240 -5068 291 -5030
rect 240 -1518 291 -1480
rect 240 -8121 291 -8083
rect 240 -3719 291 -3681
rect 240 -1873 291 -1835
rect 240 -8405 291 -8367
rect 240 -6062 291 -6024
rect 240 -1376 291 -1338
rect 240 -8618 291 -8580
rect 240 -1589 291 -1551
rect 240 -1447 291 -1409
rect 240 -2086 291 -2048
rect 240 -7127 291 -7089
rect 240 -1163 291 -1125
rect 240 -4003 291 -3965
rect 240 -4997 291 -4959
rect 240 -7340 291 -7302
rect 240 -1731 291 -1693
rect 240 -2512 291 -2474
rect 240 -4926 291 -4888
rect 240 -3506 291 -3468
rect 240 -1660 291 -1622
rect 240 -3080 291 -3042
rect 240 -8050 291 -8012
rect 240 -3151 291 -3113
rect 240 -4358 291 -4320
rect 240 -7837 291 -7799
rect 240 -2796 291 -2758
rect 240 -6133 291 -6095
rect 240 -1802 291 -1764
rect 157 -3435 208 -3397
rect 157 -8334 208 -8296
rect 157 -6772 208 -6734
rect 157 -2157 208 -2119
rect 157 -1305 208 -1267
rect 157 -3648 208 -3610
rect 157 -2725 208 -2687
rect 157 -3222 208 -3184
rect 157 -7766 208 -7728
rect 157 -5636 208 -5598
rect 157 -7624 208 -7586
rect 157 -7908 208 -7870
rect 157 -1234 208 -1196
rect 157 -5210 208 -5172
rect 157 -2228 208 -2190
rect 157 -5707 208 -5669
rect 157 -3577 208 -3539
rect 157 -6346 208 -6308
rect 157 -2867 208 -2829
rect 157 -6630 208 -6592
rect 157 -6417 208 -6379
rect 157 -6701 208 -6663
rect 157 -4074 208 -4036
rect 157 -8263 208 -8225
rect 157 -7979 208 -7941
rect 157 -1944 208 -1906
rect 157 -6488 208 -6450
rect 157 -5565 208 -5527
rect 157 -5494 208 -5456
rect 157 -3364 208 -3326
rect 157 -2015 208 -1977
rect 157 -5352 208 -5314
rect 157 -1518 208 -1480
rect 157 -8121 208 -8083
rect 157 -7269 208 -7231
rect 157 -1873 208 -1835
rect 157 -5423 208 -5385
rect 157 -1376 208 -1338
rect 157 -8618 208 -8580
rect 157 -1589 208 -1551
rect 157 -1447 208 -1409
rect 157 -2086 208 -2048
rect 157 -1163 208 -1125
rect 157 -3293 208 -3255
rect 157 -4003 208 -3965
rect 157 -7340 208 -7302
rect 157 -1731 208 -1693
rect 157 -3506 208 -3468
rect 157 -4145 208 -4107
rect 157 -1660 208 -1622
rect 157 -8050 208 -8012
rect 157 -8689 208 -8651
rect 157 -7837 208 -7799
rect 157 -6559 208 -6521
rect 157 -4216 208 -4178
rect 157 -2654 208 -2616
rect 157 -5281 208 -5243
rect 157 -2796 208 -2758
rect 157 -8192 208 -8154
rect 157 -7695 208 -7657
rect 157 -1802 208 -1764
rect -9 -3435 42 -3397
rect -9 -5920 42 -5882
rect -9 -6772 42 -6734
rect -9 -8334 42 -8296
rect -9 -2157 42 -2119
rect -9 -1305 42 -1267
rect -9 -3648 42 -3610
rect -9 -3222 42 -3184
rect -9 -5849 42 -5811
rect -9 -6204 42 -6166
rect -9 -7766 42 -7728
rect -9 -7624 42 -7586
rect -9 -8192 42 -8154
rect -9 -8476 42 -8438
rect -9 -7908 42 -7870
rect -9 -1234 42 -1196
rect -9 -2228 42 -2190
rect -9 -3577 42 -3539
rect -9 -6275 42 -6237
rect -9 -6346 42 -6308
rect -9 -6630 42 -6592
rect -9 -2938 42 -2900
rect -9 -6417 42 -6379
rect -9 -6701 42 -6663
rect -9 -3861 42 -3823
rect -9 -8263 42 -8225
rect -9 -5778 42 -5740
rect -9 -1944 42 -1906
rect -9 -7979 42 -7941
rect -9 -6488 42 -6450
rect -9 -3790 42 -3752
rect -9 -8547 42 -8509
rect -9 -7553 42 -7515
rect -9 -3364 42 -3326
rect -9 -2015 42 -1977
rect -9 -1518 42 -1480
rect -9 -5991 42 -5953
rect -9 -8121 42 -8083
rect -9 -3009 42 -2971
rect -9 -3932 42 -3894
rect -9 -3719 42 -3681
rect -9 -1873 42 -1835
rect -9 -8405 42 -8367
rect -9 -6062 42 -6024
rect -9 -1376 42 -1338
rect -9 -1589 42 -1551
rect -9 -1447 42 -1409
rect -9 -2086 42 -2048
rect -9 -7482 42 -7444
rect -9 -1163 42 -1125
rect -9 -3293 42 -3255
rect -9 -1731 42 -1693
rect -9 -3506 42 -3468
rect -9 -1660 42 -1622
rect -9 -3080 42 -3042
rect -9 -8050 42 -8012
rect -9 -3151 42 -3113
rect -9 -7837 42 -7799
rect -9 -6559 42 -6521
rect -9 -6133 42 -6095
rect -9 -7411 42 -7373
rect -9 -7695 42 -7657
rect -9 -1802 42 -1764
<< ndcontact >>
rect 91 -1188 108 -1171
rect 838 -1188 855 -1171
rect 589 -1188 606 -1171
rect 340 -1188 357 -1171
rect 91 -1330 108 -1313
rect 838 -1330 855 -1313
rect 589 -1330 606 -1313
rect 340 -1330 357 -1313
rect 91 -1472 108 -1455
rect 838 -1472 855 -1455
rect 589 -1472 606 -1455
rect 340 -1472 357 -1455
rect 91 -1614 108 -1597
rect 838 -1614 855 -1597
rect 589 -1614 606 -1597
rect 340 -1614 357 -1597
rect 91 -1756 108 -1739
rect 838 -1756 855 -1739
rect 589 -1756 606 -1739
rect 340 -1756 357 -1739
rect 91 -1898 108 -1881
rect 838 -1898 855 -1881
rect 589 -1898 606 -1881
rect 340 -1898 357 -1881
rect 91 -2040 108 -2023
rect 838 -2040 855 -2023
rect 589 -2040 606 -2023
rect 340 -2040 357 -2023
rect 91 -2182 108 -2165
rect 838 -2182 855 -2165
rect 589 -2182 606 -2165
rect 340 -2182 357 -2165
rect 838 -2324 855 -2307
rect 589 -2324 606 -2307
rect 838 -2466 855 -2449
rect 589 -2466 606 -2449
rect 340 -2466 357 -2449
rect 91 -2608 108 -2591
rect 838 -2608 855 -2591
rect 589 -2608 606 -2591
rect 340 -2608 357 -2591
rect 91 -2750 108 -2733
rect 838 -2750 855 -2733
rect 589 -2750 606 -2733
rect 340 -2750 357 -2733
rect 91 -2892 108 -2875
rect 838 -2892 855 -2875
rect 589 -2892 606 -2875
rect 340 -2892 357 -2875
rect 91 -3034 108 -3017
rect 838 -3034 855 -3017
rect 589 -3034 606 -3017
rect 340 -3034 357 -3017
rect 91 -3176 108 -3159
rect 838 -3176 855 -3159
rect 589 -3176 606 -3159
rect 340 -3176 357 -3159
rect 91 -3318 108 -3301
rect 838 -3318 855 -3301
rect 589 -3318 606 -3301
rect 340 -3318 357 -3301
rect 91 -3460 108 -3443
rect 838 -3460 855 -3443
rect 589 -3460 606 -3443
rect 340 -3460 357 -3443
rect 91 -3602 108 -3585
rect 838 -3602 855 -3585
rect 589 -3602 606 -3585
rect 340 -3602 357 -3585
rect 91 -3744 108 -3727
rect 838 -3744 855 -3727
rect 589 -3744 606 -3727
rect 340 -3744 357 -3727
rect 91 -3886 108 -3869
rect 838 -3886 855 -3869
rect 589 -3886 606 -3869
rect 340 -3886 357 -3869
rect 91 -4028 108 -4011
rect 838 -4028 855 -4011
rect 589 -4028 606 -4011
rect 340 -4028 357 -4011
rect 91 -4170 108 -4153
rect 838 -4170 855 -4153
rect 589 -4170 606 -4153
rect 340 -4170 357 -4153
rect 838 -4312 855 -4295
rect 589 -4312 606 -4295
rect 340 -4312 357 -4295
rect 838 -4454 855 -4437
rect 589 -4454 606 -4437
rect 340 -4454 357 -4437
rect 838 -4596 855 -4579
rect 589 -4596 606 -4579
rect 838 -4738 855 -4721
rect 589 -4738 606 -4721
rect 340 -4738 357 -4721
rect 838 -4880 855 -4863
rect 589 -4880 606 -4863
rect 340 -4880 357 -4863
rect 838 -5022 855 -5005
rect 589 -5022 606 -5005
rect 340 -5022 357 -5005
rect 91 -5164 108 -5147
rect 838 -5164 855 -5147
rect 589 -5164 606 -5147
rect 340 -5164 357 -5147
rect 91 -5306 108 -5289
rect 838 -5306 855 -5289
rect 589 -5306 606 -5289
rect 340 -5306 357 -5289
rect 91 -5448 108 -5431
rect 838 -5448 855 -5431
rect 589 -5448 606 -5431
rect 340 -5448 357 -5431
rect 91 -5590 108 -5573
rect 838 -5590 855 -5573
rect 589 -5590 606 -5573
rect 340 -5590 357 -5573
rect 91 -5732 108 -5715
rect 838 -5732 855 -5715
rect 589 -5732 606 -5715
rect 340 -5732 357 -5715
rect 91 -5874 108 -5857
rect 838 -5874 855 -5857
rect 589 -5874 606 -5857
rect 340 -5874 357 -5857
rect 91 -6016 108 -5999
rect 838 -6016 855 -5999
rect 589 -6016 606 -5999
rect 340 -6016 357 -5999
rect 91 -6158 108 -6141
rect 838 -6158 855 -6141
rect 589 -6158 606 -6141
rect 340 -6158 357 -6141
rect 91 -6300 108 -6283
rect 838 -6300 855 -6283
rect 589 -6300 606 -6283
rect 340 -6300 357 -6283
rect 91 -6442 108 -6425
rect 838 -6442 855 -6425
rect 589 -6442 606 -6425
rect 340 -6442 357 -6425
rect 91 -6584 108 -6567
rect 838 -6584 855 -6567
rect 589 -6584 606 -6567
rect 340 -6584 357 -6567
rect 91 -6726 108 -6709
rect 838 -6726 855 -6709
rect 589 -6726 606 -6709
rect 340 -6726 357 -6709
rect 838 -6868 855 -6851
rect 838 -7010 855 -6993
rect 589 -7010 606 -6993
rect 340 -7010 357 -6993
rect 838 -7152 855 -7135
rect 589 -7152 606 -7135
rect 340 -7152 357 -7135
rect 91 -7294 108 -7277
rect 838 -7294 855 -7277
rect 589 -7294 606 -7277
rect 340 -7294 357 -7277
rect 91 -7436 108 -7419
rect 589 -7436 606 -7419
rect 340 -7436 357 -7419
rect 91 -7578 108 -7561
rect 838 -7578 855 -7561
rect 589 -7578 606 -7561
rect 340 -7578 357 -7561
rect 91 -7720 108 -7703
rect 838 -7720 855 -7703
rect 589 -7720 606 -7703
rect 340 -7720 357 -7703
rect 91 -7862 108 -7845
rect 838 -7862 855 -7845
rect 589 -7862 606 -7845
rect 340 -7862 357 -7845
rect 91 -8004 108 -7987
rect 838 -8004 855 -7987
rect 589 -8004 606 -7987
rect 340 -8004 357 -7987
rect 91 -8146 108 -8129
rect 838 -8146 855 -8129
rect 589 -8146 606 -8129
rect 340 -8146 357 -8129
rect 91 -8288 108 -8271
rect 838 -8288 855 -8271
rect 589 -8288 606 -8271
rect 340 -8288 357 -8271
rect 91 -8430 108 -8413
rect 589 -8430 606 -8413
rect 340 -8430 357 -8413
rect 91 -8572 108 -8555
rect 838 -8572 855 -8555
rect 589 -8572 606 -8555
rect 340 -8572 357 -8555
rect 91 -8714 108 -8697
rect 838 -8714 855 -8697
rect 589 -8714 606 -8697
rect 340 -8714 357 -8697
rect 838 -8856 855 -8839
rect 589 -8856 606 -8839
rect 340 -8856 357 -8839
rect 838 -8998 855 -8981
rect 589 -8998 606 -8981
rect 672 -1117 689 -1100
rect 921 -1117 938 -1100
rect 506 -1117 523 -1100
rect 755 -1117 772 -1100
rect 174 -1117 191 -1100
rect 423 -1117 440 -1100
rect 8 -1117 25 -1100
rect 257 -1117 274 -1100
rect 672 -1259 689 -1242
rect 921 -1259 938 -1242
rect 506 -1259 523 -1242
rect 755 -1259 772 -1242
rect 174 -1259 191 -1242
rect 423 -1259 440 -1242
rect 8 -1259 25 -1242
rect 257 -1259 274 -1242
rect 672 -1401 689 -1384
rect 921 -1401 938 -1384
rect 506 -1401 523 -1384
rect 755 -1401 772 -1384
rect 174 -1401 191 -1384
rect 423 -1401 440 -1384
rect 8 -1401 25 -1384
rect 257 -1401 274 -1384
rect 672 -1543 689 -1526
rect 921 -1543 938 -1526
rect 506 -1543 523 -1526
rect 755 -1543 772 -1526
rect 174 -1543 191 -1526
rect 423 -1543 440 -1526
rect 8 -1543 25 -1526
rect 257 -1543 274 -1526
rect 672 -1685 689 -1668
rect 921 -1685 938 -1668
rect 506 -1685 523 -1668
rect 755 -1685 772 -1668
rect 174 -1685 191 -1668
rect 423 -1685 440 -1668
rect 8 -1685 25 -1668
rect 257 -1685 274 -1668
rect 672 -1827 689 -1810
rect 921 -1827 938 -1810
rect 506 -1827 523 -1810
rect 755 -1827 772 -1810
rect 174 -1827 191 -1810
rect 423 -1827 440 -1810
rect 8 -1827 25 -1810
rect 257 -1827 274 -1810
rect 672 -1969 689 -1952
rect 921 -1969 938 -1952
rect 506 -1969 523 -1952
rect 755 -1969 772 -1952
rect 174 -1969 191 -1952
rect 423 -1969 440 -1952
rect 8 -1969 25 -1952
rect 257 -1969 274 -1952
rect 672 -2111 689 -2094
rect 921 -2111 938 -2094
rect 506 -2111 523 -2094
rect 755 -2111 772 -2094
rect 174 -2111 191 -2094
rect 423 -2111 440 -2094
rect 8 -2111 25 -2094
rect 257 -2111 274 -2094
rect 672 -2253 689 -2236
rect 921 -2253 938 -2236
rect 506 -2253 523 -2236
rect 755 -2253 772 -2236
rect 174 -2253 191 -2236
rect 423 -2253 440 -2236
rect 8 -2253 25 -2236
rect 257 -2253 274 -2236
rect 672 -2395 689 -2378
rect 921 -2395 938 -2378
rect 506 -2395 523 -2378
rect 755 -2395 772 -2378
rect 423 -2395 440 -2378
rect 672 -2537 689 -2520
rect 921 -2537 938 -2520
rect 506 -2537 523 -2520
rect 755 -2537 772 -2520
rect 423 -2537 440 -2520
rect 257 -2537 274 -2520
rect 672 -2679 689 -2662
rect 921 -2679 938 -2662
rect 506 -2679 523 -2662
rect 755 -2679 772 -2662
rect 174 -2679 191 -2662
rect 423 -2679 440 -2662
rect 672 -2821 689 -2804
rect 921 -2821 938 -2804
rect 506 -2821 523 -2804
rect 755 -2821 772 -2804
rect 174 -2821 191 -2804
rect 423 -2821 440 -2804
rect 257 -2821 274 -2804
rect 672 -2963 689 -2946
rect 921 -2963 938 -2946
rect 506 -2963 523 -2946
rect 755 -2963 772 -2946
rect 423 -2963 440 -2946
rect 8 -2963 25 -2946
rect 672 -3105 689 -3088
rect 921 -3105 938 -3088
rect 506 -3105 523 -3088
rect 755 -3105 772 -3088
rect 423 -3105 440 -3088
rect 8 -3105 25 -3088
rect 257 -3105 274 -3088
rect 672 -3247 689 -3230
rect 921 -3247 938 -3230
rect 506 -3247 523 -3230
rect 755 -3247 772 -3230
rect 174 -3247 191 -3230
rect 423 -3247 440 -3230
rect 8 -3247 25 -3230
rect 672 -3389 689 -3372
rect 921 -3389 938 -3372
rect 506 -3389 523 -3372
rect 755 -3389 772 -3372
rect 174 -3389 191 -3372
rect 423 -3389 440 -3372
rect 8 -3389 25 -3372
rect 257 -3389 274 -3372
rect 672 -3531 689 -3514
rect 921 -3531 938 -3514
rect 506 -3531 523 -3514
rect 755 -3531 772 -3514
rect 174 -3531 191 -3514
rect 423 -3531 440 -3514
rect 8 -3531 25 -3514
rect 257 -3531 274 -3514
rect 672 -3673 689 -3656
rect 921 -3673 938 -3656
rect 506 -3673 523 -3656
rect 755 -3673 772 -3656
rect 174 -3673 191 -3656
rect 423 -3673 440 -3656
rect 8 -3673 25 -3656
rect 257 -3673 274 -3656
rect 672 -3815 689 -3798
rect 921 -3815 938 -3798
rect 506 -3815 523 -3798
rect 755 -3815 772 -3798
rect 423 -3815 440 -3798
rect 8 -3815 25 -3798
rect 257 -3815 274 -3798
rect 672 -3957 689 -3940
rect 921 -3957 938 -3940
rect 506 -3957 523 -3940
rect 755 -3957 772 -3940
rect 174 -3957 191 -3940
rect 423 -3957 440 -3940
rect 8 -3957 25 -3940
rect 257 -3957 274 -3940
rect 672 -4099 689 -4082
rect 921 -4099 938 -4082
rect 506 -4099 523 -4082
rect 755 -4099 772 -4082
rect 174 -4099 191 -4082
rect 423 -4099 440 -4082
rect 257 -4099 274 -4082
rect 672 -4241 689 -4224
rect 921 -4241 938 -4224
rect 506 -4241 523 -4224
rect 755 -4241 772 -4224
rect 174 -4241 191 -4224
rect 423 -4241 440 -4224
rect 257 -4241 274 -4224
rect 672 -4383 689 -4366
rect 921 -4383 938 -4366
rect 506 -4383 523 -4366
rect 755 -4383 772 -4366
rect 423 -4383 440 -4366
rect 257 -4383 274 -4366
rect 672 -4525 689 -4508
rect 921 -4525 938 -4508
rect 506 -4525 523 -4508
rect 755 -4525 772 -4508
rect 672 -4667 689 -4650
rect 921 -4667 938 -4650
rect 506 -4667 523 -4650
rect 755 -4667 772 -4650
rect 672 -4809 689 -4792
rect 921 -4809 938 -4792
rect 506 -4809 523 -4792
rect 755 -4809 772 -4792
rect 423 -4809 440 -4792
rect 672 -4951 689 -4934
rect 921 -4951 938 -4934
rect 506 -4951 523 -4934
rect 755 -4951 772 -4934
rect 257 -4951 274 -4934
rect 672 -5093 689 -5076
rect 921 -5093 938 -5076
rect 506 -5093 523 -5076
rect 755 -5093 772 -5076
rect 423 -5093 440 -5076
rect 257 -5093 274 -5076
rect 672 -5235 689 -5218
rect 921 -5235 938 -5218
rect 506 -5235 523 -5218
rect 755 -5235 772 -5218
rect 174 -5235 191 -5218
rect 672 -5377 689 -5360
rect 921 -5377 938 -5360
rect 506 -5377 523 -5360
rect 755 -5377 772 -5360
rect 174 -5377 191 -5360
rect 423 -5377 440 -5360
rect 672 -5519 689 -5502
rect 921 -5519 938 -5502
rect 506 -5519 523 -5502
rect 755 -5519 772 -5502
rect 174 -5519 191 -5502
rect 257 -5519 274 -5502
rect 672 -5661 689 -5644
rect 921 -5661 938 -5644
rect 506 -5661 523 -5644
rect 755 -5661 772 -5644
rect 174 -5661 191 -5644
rect 423 -5661 440 -5644
rect 257 -5661 274 -5644
rect 672 -5803 689 -5786
rect 921 -5803 938 -5786
rect 506 -5803 523 -5786
rect 755 -5803 772 -5786
rect 8 -5803 25 -5786
rect 672 -5945 689 -5928
rect 921 -5945 938 -5928
rect 506 -5945 523 -5928
rect 755 -5945 772 -5928
rect 423 -5945 440 -5928
rect 8 -5945 25 -5928
rect 672 -6087 689 -6070
rect 921 -6087 938 -6070
rect 506 -6087 523 -6070
rect 755 -6087 772 -6070
rect 8 -6087 25 -6070
rect 257 -6087 274 -6070
rect 672 -6229 689 -6212
rect 921 -6229 938 -6212
rect 506 -6229 523 -6212
rect 755 -6229 772 -6212
rect 423 -6229 440 -6212
rect 8 -6229 25 -6212
rect 257 -6229 274 -6212
rect 672 -6371 689 -6354
rect 921 -6371 938 -6354
rect 506 -6371 523 -6354
rect 755 -6371 772 -6354
rect 174 -6371 191 -6354
rect 8 -6371 25 -6354
rect 672 -6513 689 -6496
rect 921 -6513 938 -6496
rect 506 -6513 523 -6496
rect 755 -6513 772 -6496
rect 174 -6513 191 -6496
rect 423 -6513 440 -6496
rect 8 -6513 25 -6496
rect 672 -6655 689 -6638
rect 921 -6655 938 -6638
rect 506 -6655 523 -6638
rect 755 -6655 772 -6638
rect 174 -6655 191 -6638
rect 8 -6655 25 -6638
rect 257 -6655 274 -6638
rect 672 -6797 689 -6780
rect 921 -6797 938 -6780
rect 755 -6797 772 -6780
rect 174 -6797 191 -6780
rect 423 -6797 440 -6780
rect 8 -6797 25 -6780
rect 257 -6797 274 -6780
rect 506 -6939 523 -6922
rect 755 -6939 772 -6922
rect 672 -7081 689 -7064
rect 921 -7081 938 -7064
rect 423 -7081 440 -7064
rect 257 -7081 274 -7064
rect 672 -7223 689 -7206
rect 921 -7223 938 -7206
rect 506 -7223 523 -7206
rect 755 -7223 772 -7206
rect 174 -7223 191 -7206
rect 423 -7223 440 -7206
rect 257 -7223 274 -7206
rect 672 -7365 689 -7348
rect 921 -7365 938 -7348
rect 755 -7365 772 -7348
rect 174 -7365 191 -7348
rect 8 -7365 25 -7348
rect 257 -7365 274 -7348
rect 506 -7507 523 -7490
rect 423 -7507 440 -7490
rect 8 -7507 25 -7490
rect 257 -7507 274 -7490
rect 672 -7649 689 -7632
rect 506 -7649 523 -7632
rect 755 -7649 772 -7632
rect 174 -7649 191 -7632
rect 423 -7649 440 -7632
rect 8 -7649 25 -7632
rect 672 -7791 689 -7774
rect 921 -7791 938 -7774
rect 506 -7791 523 -7774
rect 755 -7791 772 -7774
rect 174 -7791 191 -7774
rect 423 -7791 440 -7774
rect 8 -7791 25 -7774
rect 257 -7791 274 -7774
rect 672 -7933 689 -7916
rect 921 -7933 938 -7916
rect 506 -7933 523 -7916
rect 174 -7933 191 -7916
rect 755 -7933 772 -7916
rect 423 -7933 440 -7916
rect 8 -7933 25 -7916
rect 257 -7933 274 -7916
rect 672 -8075 689 -8058
rect 921 -8075 938 -8058
rect 506 -8075 523 -8058
rect 174 -8075 191 -8058
rect 423 -8075 440 -8058
rect 8 -8075 25 -8058
rect 257 -8075 274 -8058
rect 506 -8217 523 -8200
rect 755 -8217 772 -8200
rect 174 -8217 191 -8200
rect 423 -8217 440 -8200
rect 8 -8217 25 -8200
rect 257 -8217 274 -8200
rect 672 -8359 689 -8342
rect 755 -8359 772 -8342
rect 174 -8359 191 -8342
rect 423 -8359 440 -8342
rect 8 -8359 25 -8342
rect 257 -8359 274 -8342
rect 506 -8501 523 -8484
rect 423 -8501 440 -8484
rect 8 -8501 25 -8484
rect 672 -8643 689 -8626
rect 921 -8643 938 -8626
rect 506 -8643 523 -8626
rect 755 -8643 772 -8626
rect 174 -8643 191 -8626
rect 257 -8643 274 -8626
rect 672 -8785 689 -8768
rect 921 -8785 938 -8768
rect 506 -8785 523 -8768
rect 423 -8785 440 -8768
rect 257 -8785 274 -8768
rect 672 -8927 689 -8910
rect 921 -8927 938 -8910
rect 506 -8927 523 -8910
rect 755 -8927 772 -8910
rect 423 -8927 440 -8910
rect 755 -9069 772 -9052
<< end >>