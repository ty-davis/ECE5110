* NGSPICE file created from tristate.ext - technology: sky130A

*.subckt tristate VDD GND A Y EN ~EN
X0 a_174_130# A GND GND sky130_fd_pr__nfet_01v8 ad=0.0525 pd=0.71 as=0.18 ps=1.72 w=0.5 l=0.15
X1 a_174_630# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 Y ~EN a_174_630# VDD sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.72 as=0.195 ps=1.39 w=1 l=0.15
X3 Y EN a_174_130# GND sky130_fd_pr__nfet_01v8 ad=0.18 pd=1.72 as=0.0525 ps=0.71 w=0.5 l=0.15
*.ends

