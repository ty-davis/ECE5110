magic
tech sky130A
timestamp 1744679307
<< nwell >>
rect -27 120 973 300
<< nmos >>
<< pmos >>
<< ndiff >>
rect 830 -9148 863 -9115
rect 489 -9148 581 -9115
rect 365 -9148 457 -9115
rect 332 -9148 365 -9115
rect -9 -9148 83 -9115
rect 83 -9148 116 -9115
rect 116 -9148 208 -9115
rect 614 -9148 706 -9115
rect 581 -9148 614 -9115
rect 738 -9148 830 -9115
rect 240 -9148 332 -9115
rect 863 -9148 955 -9115
rect 830 -9290 863 -9257
rect 489 -9290 581 -9257
rect 365 -9290 457 -9257
rect 332 -9290 365 -9257
rect -9 -9290 83 -9257
rect 83 -9290 116 -9257
rect 116 -9290 208 -9257
rect 614 -9290 706 -9257
rect 581 -9290 614 -9257
rect 738 -9290 830 -9257
rect 240 -9290 332 -9257
rect 863 -9290 955 -9257
rect 830 -9432 863 -9399
rect 489 -9432 581 -9399
rect 365 -9432 457 -9399
rect 332 -9432 365 -9399
rect -9 -9432 83 -9399
rect 83 -9432 116 -9399
rect 116 -9432 208 -9399
rect 614 -9432 706 -9399
rect 581 -9432 614 -9399
rect 738 -9432 830 -9399
rect 240 -9432 332 -9399
rect 863 -9432 955 -9399
rect 830 -9574 863 -9541
rect 489 -9574 581 -9541
rect 365 -9574 457 -9541
rect 332 -9574 365 -9541
rect -9 -9574 83 -9541
rect 83 -9574 116 -9541
rect 116 -9574 208 -9541
rect 614 -9574 706 -9541
rect 581 -9574 614 -9541
rect 738 -9574 830 -9541
rect 240 -9574 332 -9541
rect 863 -9574 955 -9541
rect 830 -9716 863 -9683
rect 489 -9716 581 -9683
rect 365 -9716 457 -9683
rect 332 -9716 365 -9683
rect -9 -9716 83 -9683
rect 83 -9716 116 -9683
rect 116 -9716 208 -9683
rect 614 -9716 706 -9683
rect 581 -9716 614 -9683
rect 738 -9716 830 -9683
rect 240 -9716 332 -9683
rect 863 -9716 955 -9683
rect 830 -9858 863 -9825
rect 489 -9858 581 -9825
rect 365 -9858 457 -9825
rect 332 -9858 365 -9825
rect -9 -9858 83 -9825
rect 83 -9858 116 -9825
rect 116 -9858 208 -9825
rect 614 -9858 706 -9825
rect 581 -9858 614 -9825
rect 738 -9858 830 -9825
rect 240 -9858 332 -9825
rect 863 -9858 955 -9825
rect 830 -10000 863 -9967
rect 489 -10000 581 -9967
rect 365 -10000 457 -9967
rect 332 -10000 365 -9967
rect -9 -10000 83 -9967
rect 83 -10000 116 -9967
rect 116 -10000 208 -9967
rect 614 -10000 706 -9967
rect 581 -10000 614 -9967
rect 738 -10000 830 -9967
rect 240 -10000 332 -9967
rect 863 -10000 955 -9967
rect 830 -10142 863 -10109
rect 489 -10142 581 -10109
rect 365 -10142 457 -10109
rect 332 -10142 365 -10109
rect -9 -10142 83 -10109
rect 83 -10142 116 -10109
rect 116 -10142 208 -10109
rect 614 -10142 706 -10109
rect 581 -10142 614 -10109
rect 738 -10142 830 -10109
rect 240 -10142 332 -10109
rect 863 -10142 955 -10109
rect 830 -10284 863 -10251
rect 489 -10284 581 -10251
rect 365 -10284 457 -10251
rect 332 -10284 365 -10251
rect -9 -10284 83 -10251
rect 83 -10284 116 -10251
rect 116 -10284 208 -10251
rect 614 -10284 706 -10251
rect 581 -10284 614 -10251
rect 738 -10284 830 -10251
rect 240 -10284 332 -10251
rect 863 -10284 955 -10251
rect 830 -10426 863 -10393
rect 489 -10426 581 -10393
rect 365 -10426 457 -10393
rect 332 -10426 365 -10393
rect -9 -10426 83 -10393
rect 83 -10426 116 -10393
rect 116 -10426 208 -10393
rect 614 -10426 706 -10393
rect 581 -10426 614 -10393
rect 738 -10426 830 -10393
rect 240 -10426 332 -10393
rect 863 -10426 955 -10393
rect 830 -10568 863 -10535
rect 489 -10568 581 -10535
rect 365 -10568 457 -10535
rect 332 -10568 365 -10535
rect -9 -10568 83 -10535
rect 83 -10568 116 -10535
rect 116 -10568 208 -10535
rect 614 -10568 706 -10535
rect 581 -10568 614 -10535
rect 738 -10568 830 -10535
rect 240 -10568 332 -10535
rect 863 -10568 955 -10535
rect 830 -10710 863 -10677
rect 489 -10710 581 -10677
rect 365 -10710 457 -10677
rect 332 -10710 365 -10677
rect -9 -10710 83 -10677
rect 83 -10710 116 -10677
rect 116 -10710 208 -10677
rect 614 -10710 706 -10677
rect 581 -10710 614 -10677
rect 738 -10710 830 -10677
rect 240 -10710 332 -10677
rect 863 -10710 955 -10677
rect 830 -10852 863 -10819
rect 489 -10852 581 -10819
rect 365 -10852 457 -10819
rect 332 -10852 365 -10819
rect -9 -10852 83 -10819
rect 83 -10852 116 -10819
rect 116 -10852 208 -10819
rect 614 -10852 706 -10819
rect 581 -10852 614 -10819
rect 738 -10852 830 -10819
rect 240 -10852 332 -10819
rect 863 -10852 955 -10819
rect 830 -10994 863 -10961
rect 489 -10994 581 -10961
rect 365 -10994 457 -10961
rect 332 -10994 365 -10961
rect -9 -10994 83 -10961
rect 83 -10994 116 -10961
rect 116 -10994 208 -10961
rect 614 -10994 706 -10961
rect 581 -10994 614 -10961
rect 738 -10994 830 -10961
rect 240 -10994 332 -10961
rect 863 -10994 955 -10961
rect 830 -11136 863 -11103
rect 489 -11136 581 -11103
rect 365 -11136 457 -11103
rect 332 -11136 365 -11103
rect -9 -11136 83 -11103
rect 83 -11136 116 -11103
rect 116 -11136 208 -11103
rect 614 -11136 706 -11103
rect 581 -11136 614 -11103
rect 738 -11136 830 -11103
rect 240 -11136 332 -11103
rect 863 -11136 955 -11103
rect 830 -11278 863 -11245
rect 489 -11278 581 -11245
rect 365 -11278 457 -11245
rect 332 -11278 365 -11245
rect -9 -11278 83 -11245
rect 83 -11278 116 -11245
rect 116 -11278 208 -11245
rect 614 -11278 706 -11245
rect 581 -11278 614 -11245
rect 738 -11278 830 -11245
rect 240 -11278 332 -11245
rect 863 -11278 955 -11245
rect 830 -11420 863 -11387
rect 489 -11420 581 -11387
rect 365 -11420 457 -11387
rect 332 -11420 365 -11387
rect -9 -11420 83 -11387
rect 83 -11420 116 -11387
rect 116 -11420 208 -11387
rect 614 -11420 706 -11387
rect 581 -11420 614 -11387
rect 738 -11420 830 -11387
rect 240 -11420 332 -11387
rect 863 -11420 955 -11387
rect 830 -11562 863 -11529
rect 489 -11562 581 -11529
rect 365 -11562 457 -11529
rect 332 -11562 365 -11529
rect -9 -11562 83 -11529
rect 83 -11562 116 -11529
rect 116 -11562 208 -11529
rect 614 -11562 706 -11529
rect 581 -11562 614 -11529
rect 738 -11562 830 -11529
rect 240 -11562 332 -11529
rect 863 -11562 955 -11529
rect 830 -11704 863 -11671
rect 489 -11704 581 -11671
rect 365 -11704 457 -11671
rect 332 -11704 365 -11671
rect -9 -11704 83 -11671
rect 83 -11704 116 -11671
rect 116 -11704 208 -11671
rect 614 -11704 706 -11671
rect 581 -11704 614 -11671
rect 738 -11704 830 -11671
rect 240 -11704 332 -11671
rect 863 -11704 955 -11671
rect 830 -11846 863 -11813
rect 489 -11846 581 -11813
rect 365 -11846 457 -11813
rect 332 -11846 365 -11813
rect -9 -11846 83 -11813
rect 83 -11846 116 -11813
rect 116 -11846 208 -11813
rect 614 -11846 706 -11813
rect 581 -11846 614 -11813
rect 738 -11846 830 -11813
rect 240 -11846 332 -11813
rect 863 -11846 955 -11813
rect 830 -11988 863 -11955
rect 489 -11988 581 -11955
rect 365 -11988 457 -11955
rect 332 -11988 365 -11955
rect -9 -11988 83 -11955
rect 83 -11988 116 -11955
rect 116 -11988 208 -11955
rect 614 -11988 706 -11955
rect 581 -11988 614 -11955
rect 738 -11988 830 -11955
rect 240 -11988 332 -11955
rect 863 -11988 955 -11955
rect 830 -12130 863 -12097
rect 489 -12130 581 -12097
rect 365 -12130 457 -12097
rect 332 -12130 365 -12097
rect -9 -12130 83 -12097
rect 83 -12130 116 -12097
rect 116 -12130 208 -12097
rect 614 -12130 706 -12097
rect 581 -12130 614 -12097
rect 738 -12130 830 -12097
rect 240 -12130 332 -12097
rect 863 -12130 955 -12097
rect 830 -12272 863 -12239
rect 489 -12272 581 -12239
rect 365 -12272 457 -12239
rect 332 -12272 365 -12239
rect -9 -12272 83 -12239
rect 83 -12272 116 -12239
rect 116 -12272 208 -12239
rect 614 -12272 706 -12239
rect 581 -12272 614 -12239
rect 738 -12272 830 -12239
rect 240 -12272 332 -12239
rect 863 -12272 955 -12239
rect 830 -12414 863 -12381
rect 489 -12414 581 -12381
rect 365 -12414 457 -12381
rect 332 -12414 365 -12381
rect -9 -12414 83 -12381
rect 83 -12414 116 -12381
rect 116 -12414 208 -12381
rect 614 -12414 706 -12381
rect 581 -12414 614 -12381
rect 738 -12414 830 -12381
rect 240 -12414 332 -12381
rect 863 -12414 955 -12381
rect 830 -12556 863 -12523
rect 489 -12556 581 -12523
rect 365 -12556 457 -12523
rect 332 -12556 365 -12523
rect -9 -12556 83 -12523
rect 83 -12556 116 -12523
rect 116 -12556 208 -12523
rect 614 -12556 706 -12523
rect 581 -12556 614 -12523
rect 738 -12556 830 -12523
rect 240 -12556 332 -12523
rect 863 -12556 955 -12523
rect 830 -12698 863 -12665
rect 489 -12698 581 -12665
rect 365 -12698 457 -12665
rect 332 -12698 365 -12665
rect -9 -12698 83 -12665
rect 83 -12698 116 -12665
rect 116 -12698 208 -12665
rect 614 -12698 706 -12665
rect 581 -12698 614 -12665
rect 738 -12698 830 -12665
rect 240 -12698 332 -12665
rect 863 -12698 955 -12665
rect 830 -12840 863 -12807
rect 489 -12840 581 -12807
rect 365 -12840 457 -12807
rect 332 -12840 365 -12807
rect -9 -12840 83 -12807
rect 83 -12840 116 -12807
rect 116 -12840 208 -12807
rect 614 -12840 706 -12807
rect 581 -12840 614 -12807
rect 738 -12840 830 -12807
rect 240 -12840 332 -12807
rect 863 -12840 955 -12807
rect 830 -12982 863 -12949
rect 489 -12982 581 -12949
rect 365 -12982 457 -12949
rect 332 -12982 365 -12949
rect -9 -12982 83 -12949
rect 83 -12982 116 -12949
rect 116 -12982 208 -12949
rect 614 -12982 706 -12949
rect 581 -12982 614 -12949
rect 738 -12982 830 -12949
rect 240 -12982 332 -12949
rect 863 -12982 955 -12949
rect 830 -13124 863 -13091
rect 489 -13124 581 -13091
rect 365 -13124 457 -13091
rect 332 -13124 365 -13091
rect -9 -13124 83 -13091
rect 83 -13124 116 -13091
rect 116 -13124 208 -13091
rect 614 -13124 706 -13091
rect 581 -13124 614 -13091
rect 738 -13124 830 -13091
rect 240 -13124 332 -13091
rect 863 -13124 955 -13091
rect 830 -13266 863 -13233
rect 489 -13266 581 -13233
rect 365 -13266 457 -13233
rect 332 -13266 365 -13233
rect -9 -13266 83 -13233
rect 83 -13266 116 -13233
rect 116 -13266 208 -13233
rect 614 -13266 706 -13233
rect 581 -13266 614 -13233
rect 738 -13266 830 -13233
rect 240 -13266 332 -13233
rect 863 -13266 955 -13233
rect 830 -13408 863 -13375
rect 489 -13408 581 -13375
rect 365 -13408 457 -13375
rect 332 -13408 365 -13375
rect -9 -13408 83 -13375
rect 83 -13408 116 -13375
rect 116 -13408 208 -13375
rect 614 -13408 706 -13375
rect 581 -13408 614 -13375
rect 738 -13408 830 -13375
rect 240 -13408 332 -13375
rect 863 -13408 955 -13375
rect 830 -13550 863 -13517
rect 489 -13550 581 -13517
rect 365 -13550 457 -13517
rect 332 -13550 365 -13517
rect -9 -13550 83 -13517
rect 83 -13550 116 -13517
rect 116 -13550 208 -13517
rect 614 -13550 706 -13517
rect 581 -13550 614 -13517
rect 738 -13550 830 -13517
rect 240 -13550 332 -13517
rect 863 -13550 955 -13517
rect 830 -13692 863 -13659
rect 489 -13692 581 -13659
rect 365 -13692 457 -13659
rect 332 -13692 365 -13659
rect -9 -13692 83 -13659
rect 83 -13692 116 -13659
rect 116 -13692 208 -13659
rect 614 -13692 706 -13659
rect 581 -13692 614 -13659
rect 738 -13692 830 -13659
rect 240 -13692 332 -13659
rect 863 -13692 955 -13659
rect 830 -13834 863 -13801
rect 489 -13834 581 -13801
rect 365 -13834 457 -13801
rect 332 -13834 365 -13801
rect -9 -13834 83 -13801
rect 83 -13834 116 -13801
rect 116 -13834 208 -13801
rect 614 -13834 706 -13801
rect 581 -13834 614 -13801
rect 738 -13834 830 -13801
rect 240 -13834 332 -13801
rect 863 -13834 955 -13801
rect 830 -13976 863 -13943
rect 489 -13976 581 -13943
rect 365 -13976 457 -13943
rect 332 -13976 365 -13943
rect -9 -13976 83 -13943
rect 83 -13976 116 -13943
rect 116 -13976 208 -13943
rect 614 -13976 706 -13943
rect 581 -13976 614 -13943
rect 738 -13976 830 -13943
rect 240 -13976 332 -13943
rect 863 -13976 955 -13943
rect 830 -14118 863 -14085
rect 489 -14118 581 -14085
rect 365 -14118 457 -14085
rect 332 -14118 365 -14085
rect -9 -14118 83 -14085
rect 83 -14118 116 -14085
rect 116 -14118 208 -14085
rect 614 -14118 706 -14085
rect 581 -14118 614 -14085
rect 738 -14118 830 -14085
rect 240 -14118 332 -14085
rect 863 -14118 955 -14085
rect 830 -14260 863 -14227
rect 489 -14260 581 -14227
rect 365 -14260 457 -14227
rect 332 -14260 365 -14227
rect -9 -14260 83 -14227
rect 83 -14260 116 -14227
rect 116 -14260 208 -14227
rect 614 -14260 706 -14227
rect 581 -14260 614 -14227
rect 738 -14260 830 -14227
rect 240 -14260 332 -14227
rect 863 -14260 955 -14227
rect 830 -14402 863 -14369
rect 489 -14402 581 -14369
rect 365 -14402 457 -14369
rect 332 -14402 365 -14369
rect -9 -14402 83 -14369
rect 83 -14402 116 -14369
rect 116 -14402 208 -14369
rect 614 -14402 706 -14369
rect 581 -14402 614 -14369
rect 738 -14402 830 -14369
rect 240 -14402 332 -14369
rect 863 -14402 955 -14369
rect 830 -14544 863 -14511
rect 489 -14544 581 -14511
rect 365 -14544 457 -14511
rect 332 -14544 365 -14511
rect -9 -14544 83 -14511
rect 83 -14544 116 -14511
rect 116 -14544 208 -14511
rect 614 -14544 706 -14511
rect 581 -14544 614 -14511
rect 738 -14544 830 -14511
rect 240 -14544 332 -14511
rect 863 -14544 955 -14511
rect 830 -14686 863 -14653
rect 489 -14686 581 -14653
rect 365 -14686 457 -14653
rect 332 -14686 365 -14653
rect -9 -14686 83 -14653
rect 83 -14686 116 -14653
rect 116 -14686 208 -14653
rect 614 -14686 706 -14653
rect 581 -14686 614 -14653
rect 738 -14686 830 -14653
rect 240 -14686 332 -14653
rect 863 -14686 955 -14653
rect 830 -14828 863 -14795
rect 489 -14828 581 -14795
rect 365 -14828 457 -14795
rect 332 -14828 365 -14795
rect -9 -14828 83 -14795
rect 83 -14828 116 -14795
rect 116 -14828 208 -14795
rect 614 -14828 706 -14795
rect 581 -14828 614 -14795
rect 738 -14828 830 -14795
rect 240 -14828 332 -14795
rect 863 -14828 955 -14795
rect 830 -14970 863 -14937
rect 489 -14970 581 -14937
rect 365 -14970 457 -14937
rect 332 -14970 365 -14937
rect -9 -14970 83 -14937
rect 83 -14970 116 -14937
rect 116 -14970 208 -14937
rect 614 -14970 706 -14937
rect 581 -14970 614 -14937
rect 738 -14970 830 -14937
rect 240 -14970 332 -14937
rect 863 -14970 955 -14937
rect 830 -15112 863 -15079
rect 489 -15112 581 -15079
rect 365 -15112 457 -15079
rect 332 -15112 365 -15079
rect -9 -15112 83 -15079
rect 83 -15112 116 -15079
rect 116 -15112 208 -15079
rect 614 -15112 706 -15079
rect 581 -15112 614 -15079
rect 738 -15112 830 -15079
rect 240 -15112 332 -15079
rect 863 -15112 955 -15079
rect 830 -15254 863 -15221
rect 489 -15254 581 -15221
rect 365 -15254 457 -15221
rect 332 -15254 365 -15221
rect -9 -15254 83 -15221
rect 83 -15254 116 -15221
rect 116 -15254 208 -15221
rect 614 -15254 706 -15221
rect 581 -15254 614 -15221
rect 738 -15254 830 -15221
rect 240 -15254 332 -15221
rect 863 -15254 955 -15221
rect 830 -15396 863 -15363
rect 489 -15396 581 -15363
rect 365 -15396 457 -15363
rect 332 -15396 365 -15363
rect -9 -15396 83 -15363
rect 83 -15396 116 -15363
rect 116 -15396 208 -15363
rect 614 -15396 706 -15363
rect 581 -15396 614 -15363
rect 738 -15396 830 -15363
rect 240 -15396 332 -15363
rect 863 -15396 955 -15363
rect 830 -15538 863 -15505
rect 489 -15538 581 -15505
rect 365 -15538 457 -15505
rect 332 -15538 365 -15505
rect -9 -15538 83 -15505
rect 83 -15538 116 -15505
rect 116 -15538 208 -15505
rect 614 -15538 706 -15505
rect 581 -15538 614 -15505
rect 738 -15538 830 -15505
rect 240 -15538 332 -15505
rect 863 -15538 955 -15505
rect 830 -15680 863 -15647
rect 489 -15680 581 -15647
rect 365 -15680 457 -15647
rect 332 -15680 365 -15647
rect -9 -15680 83 -15647
rect 83 -15680 116 -15647
rect 116 -15680 208 -15647
rect 614 -15680 706 -15647
rect 581 -15680 614 -15647
rect 738 -15680 830 -15647
rect 240 -15680 332 -15647
rect 863 -15680 955 -15647
rect 830 -15822 863 -15789
rect 489 -15822 581 -15789
rect 365 -15822 457 -15789
rect 332 -15822 365 -15789
rect -9 -15822 83 -15789
rect 83 -15822 116 -15789
rect 116 -15822 208 -15789
rect 614 -15822 706 -15789
rect 581 -15822 614 -15789
rect 738 -15822 830 -15789
rect 240 -15822 332 -15789
rect 863 -15822 955 -15789
rect 830 -15964 863 -15931
rect 489 -15964 581 -15931
rect 365 -15964 457 -15931
rect 332 -15964 365 -15931
rect -9 -15964 83 -15931
rect 83 -15964 116 -15931
rect 116 -15964 208 -15931
rect 614 -15964 706 -15931
rect 581 -15964 614 -15931
rect 738 -15964 830 -15931
rect 240 -15964 332 -15931
rect 863 -15964 955 -15931
rect 830 -16106 863 -16073
rect 489 -16106 581 -16073
rect 365 -16106 457 -16073
rect 332 -16106 365 -16073
rect -9 -16106 83 -16073
rect 83 -16106 116 -16073
rect 116 -16106 208 -16073
rect 614 -16106 706 -16073
rect 581 -16106 614 -16073
rect 738 -16106 830 -16073
rect 240 -16106 332 -16073
rect 863 -16106 955 -16073
rect 830 -16248 863 -16215
rect 489 -16248 581 -16215
rect 365 -16248 457 -16215
rect 332 -16248 365 -16215
rect -9 -16248 83 -16215
rect 83 -16248 116 -16215
rect 116 -16248 208 -16215
rect 614 -16248 706 -16215
rect 581 -16248 614 -16215
rect 738 -16248 830 -16215
rect 240 -16248 332 -16215
rect 863 -16248 955 -16215
rect 830 -16390 863 -16357
rect 489 -16390 581 -16357
rect 365 -16390 457 -16357
rect 332 -16390 365 -16357
rect -9 -16390 83 -16357
rect 83 -16390 116 -16357
rect 116 -16390 208 -16357
rect 614 -16390 706 -16357
rect 581 -16390 614 -16357
rect 738 -16390 830 -16357
rect 240 -16390 332 -16357
rect 863 -16390 955 -16357
rect 830 -16532 863 -16499
rect 489 -16532 581 -16499
rect 365 -16532 457 -16499
rect 332 -16532 365 -16499
rect -9 -16532 83 -16499
rect 83 -16532 116 -16499
rect 116 -16532 208 -16499
rect 614 -16532 706 -16499
rect 581 -16532 614 -16499
rect 738 -16532 830 -16499
rect 240 -16532 332 -16499
rect 863 -16532 955 -16499
rect 830 -16674 863 -16641
rect 489 -16674 581 -16641
rect 365 -16674 457 -16641
rect 332 -16674 365 -16641
rect -9 -16674 83 -16641
rect 83 -16674 116 -16641
rect 116 -16674 208 -16641
rect 614 -16674 706 -16641
rect 581 -16674 614 -16641
rect 738 -16674 830 -16641
rect 240 -16674 332 -16641
rect 863 -16674 955 -16641
rect 830 -16816 863 -16783
rect 489 -16816 581 -16783
rect 365 -16816 457 -16783
rect 332 -16816 365 -16783
rect -9 -16816 83 -16783
rect 83 -16816 116 -16783
rect 116 -16816 208 -16783
rect 614 -16816 706 -16783
rect 581 -16816 614 -16783
rect 738 -16816 830 -16783
rect 240 -16816 332 -16783
rect 863 -16816 955 -16783
rect 830 -16958 863 -16925
rect 489 -16958 581 -16925
rect 365 -16958 457 -16925
rect 332 -16958 365 -16925
rect -9 -16958 83 -16925
rect 83 -16958 116 -16925
rect 116 -16958 208 -16925
rect 614 -16958 706 -16925
rect 581 -16958 614 -16925
rect 738 -16958 830 -16925
rect 240 -16958 332 -16925
rect 863 -16958 955 -16925
rect 830 -17100 863 -17067
rect 489 -17100 581 -17067
rect 365 -17100 457 -17067
rect 332 -17100 365 -17067
rect -9 -17100 83 -17067
rect 83 -17100 116 -17067
rect 116 -17100 208 -17067
rect 614 -17100 706 -17067
rect 581 -17100 614 -17067
rect 738 -17100 830 -17067
rect 240 -17100 332 -17067
rect 863 -17100 955 -17067
rect 830 -17242 863 -17209
rect 489 -17242 581 -17209
rect 365 -17242 457 -17209
rect 332 -17242 365 -17209
rect -9 -17242 83 -17209
rect 83 -17242 116 -17209
rect 116 -17242 208 -17209
rect 614 -17242 706 -17209
rect 581 -17242 614 -17209
rect 738 -17242 830 -17209
rect 240 -17242 332 -17209
rect 863 -17242 955 -17209
rect 830 -17384 863 -17351
rect 489 -17384 581 -17351
rect 365 -17384 457 -17351
rect 332 -17384 365 -17351
rect -9 -17384 83 -17351
rect 83 -17384 116 -17351
rect 116 -17384 208 -17351
rect 614 -17384 706 -17351
rect 581 -17384 614 -17351
rect 738 -17384 830 -17351
rect 240 -17384 332 -17351
rect 863 -17384 955 -17351
rect 830 -17526 863 -17493
rect 489 -17526 581 -17493
rect 365 -17526 457 -17493
rect 332 -17526 365 -17493
rect -9 -17526 83 -17493
rect 83 -17526 116 -17493
rect 116 -17526 208 -17493
rect 614 -17526 706 -17493
rect 581 -17526 614 -17493
rect 738 -17526 830 -17493
rect 240 -17526 332 -17493
rect 863 -17526 955 -17493
rect 830 -17668 863 -17635
rect 489 -17668 581 -17635
rect 365 -17668 457 -17635
rect 332 -17668 365 -17635
rect -9 -17668 83 -17635
rect 83 -17668 116 -17635
rect 116 -17668 208 -17635
rect 614 -17668 706 -17635
rect 581 -17668 614 -17635
rect 738 -17668 830 -17635
rect 240 -17668 332 -17635
rect 863 -17668 955 -17635
rect 830 -17810 863 -17777
rect 489 -17810 581 -17777
rect 365 -17810 457 -17777
rect 332 -17810 365 -17777
rect -9 -17810 83 -17777
rect 83 -17810 116 -17777
rect 116 -17810 208 -17777
rect 614 -17810 706 -17777
rect 581 -17810 614 -17777
rect 738 -17810 830 -17777
rect 240 -17810 332 -17777
rect 863 -17810 955 -17777
rect 830 -17952 863 -17919
rect 489 -17952 581 -17919
rect 365 -17952 457 -17919
rect 332 -17952 365 -17919
rect -9 -17952 83 -17919
rect 83 -17952 116 -17919
rect 116 -17952 208 -17919
rect 614 -17952 706 -17919
rect 581 -17952 614 -17919
rect 738 -17952 830 -17919
rect 240 -17952 332 -17919
rect 863 -17952 955 -17919
rect 830 -18094 863 -18061
rect 489 -18094 581 -18061
rect 365 -18094 457 -18061
rect 332 -18094 365 -18061
rect -9 -18094 83 -18061
rect 83 -18094 116 -18061
rect 116 -18094 208 -18061
rect 614 -18094 706 -18061
rect 581 -18094 614 -18061
rect 738 -18094 830 -18061
rect 240 -18094 332 -18061
rect 863 -18094 955 -18061
rect 830 -18236 863 -18203
rect 863 -18236 955 -18203
rect 830 -18378 863 -18345
rect 614 -18378 706 -18345
rect 581 -18378 614 -18345
rect 738 -18378 830 -18345
rect 863 -18378 955 -18345
rect 830 -18520 863 -18487
rect 489 -18520 581 -18487
rect 614 -18520 706 -18487
rect 581 -18520 614 -18487
rect 738 -18520 830 -18487
rect 863 -18520 955 -18487
rect 489 -18662 581 -18629
rect 830 -18662 863 -18629
rect 614 -18662 706 -18629
rect 581 -18662 614 -18629
rect 738 -18662 830 -18629
rect 863 -18662 955 -18629
rect 830 -18804 863 -18771
rect 489 -18804 581 -18771
rect 365 -18804 457 -18771
rect 332 -18804 365 -18771
rect 614 -18804 706 -18771
rect 581 -18804 614 -18771
rect 738 -18804 830 -18771
rect 863 -18804 955 -18771
rect 830 -18946 863 -18913
rect 332 -18946 365 -18913
rect 614 -18946 706 -18913
rect 365 -18946 457 -18913
rect 738 -18946 830 -18913
rect 581 -18946 614 -18913
rect 863 -18946 955 -18913
rect 830 -19088 863 -19055
rect 489 -19088 581 -19055
rect 365 -19088 457 -19055
rect 332 -19088 365 -19055
rect 614 -19088 706 -19055
rect 581 -19088 614 -19055
rect 738 -19088 830 -19055
rect 863 -19088 955 -19055
rect 489 -19230 581 -19197
rect 830 -19230 863 -19197
rect 365 -19230 457 -19197
rect 332 -19230 365 -19197
rect 614 -19230 706 -19197
rect 581 -19230 614 -19197
rect 738 -19230 830 -19197
rect 863 -19230 955 -19197
rect 830 -19372 863 -19339
rect 489 -19372 581 -19339
rect 365 -19372 457 -19339
rect 332 -19372 365 -19339
rect 614 -19372 706 -19339
rect 581 -19372 614 -19339
rect 738 -19372 830 -19339
rect 240 -19372 332 -19339
rect 863 -19372 955 -19339
rect 830 -19514 863 -19481
rect 332 -19514 365 -19481
rect 614 -19514 706 -19481
rect 581 -19514 614 -19481
rect 738 -19514 830 -19481
rect 240 -19514 332 -19481
rect 863 -19514 955 -19481
rect 830 -19656 863 -19623
rect 489 -19656 581 -19623
rect 332 -19656 365 -19623
rect 614 -19656 706 -19623
rect 581 -19656 614 -19623
rect 738 -19656 830 -19623
rect 240 -19656 332 -19623
rect 863 -19656 955 -19623
rect 489 -19798 581 -19765
rect 830 -19798 863 -19765
rect 332 -19798 365 -19765
rect 614 -19798 706 -19765
rect 581 -19798 614 -19765
rect 738 -19798 830 -19765
rect 240 -19798 332 -19765
rect 863 -19798 955 -19765
rect 830 -19940 863 -19907
rect 489 -19940 581 -19907
rect 365 -19940 457 -19907
rect 332 -19940 365 -19907
rect 614 -19940 706 -19907
rect 581 -19940 614 -19907
rect 738 -19940 830 -19907
rect 240 -19940 332 -19907
rect 863 -19940 955 -19907
rect 830 -20082 863 -20049
rect 332 -20082 365 -20049
rect 614 -20082 706 -20049
rect 365 -20082 457 -20049
rect 738 -20082 830 -20049
rect 581 -20082 614 -20049
rect 240 -20082 332 -20049
rect 863 -20082 955 -20049
rect 830 -20224 863 -20191
rect 489 -20224 581 -20191
rect 365 -20224 457 -20191
rect 332 -20224 365 -20191
rect 614 -20224 706 -20191
rect 581 -20224 614 -20191
rect 738 -20224 830 -20191
rect 240 -20224 332 -20191
rect 863 -20224 955 -20191
rect 489 -20366 581 -20333
rect 830 -20366 863 -20333
rect 365 -20366 457 -20333
rect 332 -20366 365 -20333
rect 614 -20366 706 -20333
rect 581 -20366 614 -20333
rect 738 -20366 830 -20333
rect 240 -20366 332 -20333
rect 863 -20366 955 -20333
rect 830 -20508 863 -20475
rect 489 -20508 581 -20475
rect 365 -20508 457 -20475
rect 332 -20508 365 -20475
rect 83 -20508 116 -20475
rect 116 -20508 208 -20475
rect 614 -20508 706 -20475
rect 581 -20508 614 -20475
rect 738 -20508 830 -20475
rect 240 -20508 332 -20475
rect 863 -20508 955 -20475
rect 830 -20650 863 -20617
rect 83 -20650 116 -20617
rect 116 -20650 208 -20617
rect 614 -20650 706 -20617
rect 581 -20650 614 -20617
rect 738 -20650 830 -20617
rect 863 -20650 955 -20617
rect 830 -20792 863 -20759
rect 489 -20792 581 -20759
rect 83 -20792 116 -20759
rect 116 -20792 208 -20759
rect 614 -20792 706 -20759
rect 581 -20792 614 -20759
rect 738 -20792 830 -20759
rect 863 -20792 955 -20759
rect 489 -20934 581 -20901
rect 830 -20934 863 -20901
rect 83 -20934 116 -20901
rect 116 -20934 208 -20901
rect 614 -20934 706 -20901
rect 581 -20934 614 -20901
rect 738 -20934 830 -20901
rect 863 -20934 955 -20901
rect 830 -21076 863 -21043
rect 489 -21076 581 -21043
rect 365 -21076 457 -21043
rect 332 -21076 365 -21043
rect 83 -21076 116 -21043
rect 116 -21076 208 -21043
rect 614 -21076 706 -21043
rect 581 -21076 614 -21043
rect 738 -21076 830 -21043
rect 863 -21076 955 -21043
rect 830 -21218 863 -21185
rect 332 -21218 365 -21185
rect 83 -21218 116 -21185
rect 116 -21218 208 -21185
rect 614 -21218 706 -21185
rect 365 -21218 457 -21185
rect 738 -21218 830 -21185
rect 581 -21218 614 -21185
rect 863 -21218 955 -21185
rect 830 -21360 863 -21327
rect 489 -21360 581 -21327
rect 365 -21360 457 -21327
rect 332 -21360 365 -21327
rect 83 -21360 116 -21327
rect 116 -21360 208 -21327
rect 614 -21360 706 -21327
rect 581 -21360 614 -21327
rect 738 -21360 830 -21327
rect 863 -21360 955 -21327
rect 489 -21502 581 -21469
rect 830 -21502 863 -21469
rect 365 -21502 457 -21469
rect 332 -21502 365 -21469
rect 83 -21502 116 -21469
rect 116 -21502 208 -21469
rect 614 -21502 706 -21469
rect 581 -21502 614 -21469
rect 738 -21502 830 -21469
rect 863 -21502 955 -21469
rect 830 -21644 863 -21611
rect 489 -21644 581 -21611
rect 365 -21644 457 -21611
rect 332 -21644 365 -21611
rect 83 -21644 116 -21611
rect 116 -21644 208 -21611
rect 614 -21644 706 -21611
rect 581 -21644 614 -21611
rect 738 -21644 830 -21611
rect 240 -21644 332 -21611
rect 863 -21644 955 -21611
rect 830 -21786 863 -21753
rect 332 -21786 365 -21753
rect 83 -21786 116 -21753
rect 116 -21786 208 -21753
rect 614 -21786 706 -21753
rect 581 -21786 614 -21753
rect 738 -21786 830 -21753
rect 240 -21786 332 -21753
rect 863 -21786 955 -21753
rect 830 -21928 863 -21895
rect 489 -21928 581 -21895
rect 332 -21928 365 -21895
rect 83 -21928 116 -21895
rect 116 -21928 208 -21895
rect 614 -21928 706 -21895
rect 581 -21928 614 -21895
rect 738 -21928 830 -21895
rect 240 -21928 332 -21895
rect 863 -21928 955 -21895
rect 489 -22070 581 -22037
rect 830 -22070 863 -22037
rect 332 -22070 365 -22037
rect 83 -22070 116 -22037
rect 116 -22070 208 -22037
rect 614 -22070 706 -22037
rect 581 -22070 614 -22037
rect 738 -22070 830 -22037
rect 240 -22070 332 -22037
rect 863 -22070 955 -22037
rect 830 -22212 863 -22179
rect 489 -22212 581 -22179
rect 365 -22212 457 -22179
rect 332 -22212 365 -22179
rect 83 -22212 116 -22179
rect 116 -22212 208 -22179
rect 614 -22212 706 -22179
rect 581 -22212 614 -22179
rect 738 -22212 830 -22179
rect 240 -22212 332 -22179
rect 863 -22212 955 -22179
rect 830 -22354 863 -22321
rect 332 -22354 365 -22321
rect 83 -22354 116 -22321
rect 116 -22354 208 -22321
rect 614 -22354 706 -22321
rect 365 -22354 457 -22321
rect 738 -22354 830 -22321
rect 581 -22354 614 -22321
rect 240 -22354 332 -22321
rect 863 -22354 955 -22321
rect 830 -22496 863 -22463
rect 489 -22496 581 -22463
rect 365 -22496 457 -22463
rect 332 -22496 365 -22463
rect 83 -22496 116 -22463
rect 116 -22496 208 -22463
rect 614 -22496 706 -22463
rect 581 -22496 614 -22463
rect 738 -22496 830 -22463
rect 240 -22496 332 -22463
rect 863 -22496 955 -22463
rect 489 -22638 581 -22605
rect 830 -22638 863 -22605
rect 365 -22638 457 -22605
rect 332 -22638 365 -22605
rect 83 -22638 116 -22605
rect 116 -22638 208 -22605
rect 614 -22638 706 -22605
rect 581 -22638 614 -22605
rect 738 -22638 830 -22605
rect 240 -22638 332 -22605
rect 863 -22638 955 -22605
rect 830 -22780 863 -22747
rect 489 -22780 581 -22747
rect 365 -22780 457 -22747
rect 332 -22780 365 -22747
rect -9 -22780 83 -22747
rect 83 -22780 116 -22747
rect 116 -22780 208 -22747
rect 614 -22780 706 -22747
rect 581 -22780 614 -22747
rect 738 -22780 830 -22747
rect 240 -22780 332 -22747
rect 863 -22780 955 -22747
rect 830 -22922 863 -22889
rect -9 -22922 83 -22889
rect 83 -22922 116 -22889
rect 614 -22922 706 -22889
rect 581 -22922 614 -22889
rect 738 -22922 830 -22889
rect 863 -22922 955 -22889
rect 830 -23064 863 -23031
rect 489 -23064 581 -23031
rect -9 -23064 83 -23031
rect 83 -23064 116 -23031
rect 614 -23064 706 -23031
rect 581 -23064 614 -23031
rect 738 -23064 830 -23031
rect 863 -23064 955 -23031
rect 489 -23206 581 -23173
rect 830 -23206 863 -23173
rect -9 -23206 83 -23173
rect 83 -23206 116 -23173
rect 614 -23206 706 -23173
rect 581 -23206 614 -23173
rect 738 -23206 830 -23173
rect 863 -23206 955 -23173
rect 830 -23348 863 -23315
rect 489 -23348 581 -23315
rect 365 -23348 457 -23315
rect -9 -23348 83 -23315
rect 332 -23348 365 -23315
rect 83 -23348 116 -23315
rect 614 -23348 706 -23315
rect 581 -23348 614 -23315
rect 738 -23348 830 -23315
rect 863 -23348 955 -23315
rect 830 -23490 863 -23457
rect 332 -23490 365 -23457
rect -9 -23490 83 -23457
rect 83 -23490 116 -23457
rect 614 -23490 706 -23457
rect 365 -23490 457 -23457
rect 738 -23490 830 -23457
rect 581 -23490 614 -23457
rect 863 -23490 955 -23457
rect 830 -23632 863 -23599
rect 489 -23632 581 -23599
rect 365 -23632 457 -23599
rect 332 -23632 365 -23599
rect -9 -23632 83 -23599
rect 83 -23632 116 -23599
rect 614 -23632 706 -23599
rect 581 -23632 614 -23599
rect 738 -23632 830 -23599
rect 863 -23632 955 -23599
rect 489 -23774 581 -23741
rect 830 -23774 863 -23741
rect 365 -23774 457 -23741
rect 332 -23774 365 -23741
rect -9 -23774 83 -23741
rect 83 -23774 116 -23741
rect 614 -23774 706 -23741
rect 581 -23774 614 -23741
rect 738 -23774 830 -23741
rect 863 -23774 955 -23741
rect 830 -23916 863 -23883
rect 489 -23916 581 -23883
rect 365 -23916 457 -23883
rect 332 -23916 365 -23883
rect -9 -23916 83 -23883
rect 83 -23916 116 -23883
rect 614 -23916 706 -23883
rect 581 -23916 614 -23883
rect 738 -23916 830 -23883
rect 240 -23916 332 -23883
rect 863 -23916 955 -23883
rect 830 -24058 863 -24025
rect 332 -24058 365 -24025
rect -9 -24058 83 -24025
rect 83 -24058 116 -24025
rect 614 -24058 706 -24025
rect 581 -24058 614 -24025
rect 738 -24058 830 -24025
rect 240 -24058 332 -24025
rect 863 -24058 955 -24025
rect 830 -24200 863 -24167
rect 489 -24200 581 -24167
rect 332 -24200 365 -24167
rect -9 -24200 83 -24167
rect 83 -24200 116 -24167
rect 614 -24200 706 -24167
rect 581 -24200 614 -24167
rect 738 -24200 830 -24167
rect 240 -24200 332 -24167
rect 863 -24200 955 -24167
rect 489 -24342 581 -24309
rect 830 -24342 863 -24309
rect 332 -24342 365 -24309
rect -9 -24342 83 -24309
rect 83 -24342 116 -24309
rect 614 -24342 706 -24309
rect 581 -24342 614 -24309
rect 738 -24342 830 -24309
rect 240 -24342 332 -24309
rect 863 -24342 955 -24309
rect 830 -24484 863 -24451
rect 489 -24484 581 -24451
rect 365 -24484 457 -24451
rect 332 -24484 365 -24451
rect -9 -24484 83 -24451
rect 83 -24484 116 -24451
rect 614 -24484 706 -24451
rect 581 -24484 614 -24451
rect 738 -24484 830 -24451
rect 240 -24484 332 -24451
rect 863 -24484 955 -24451
rect 830 -24626 863 -24593
rect 332 -24626 365 -24593
rect -9 -24626 83 -24593
rect 83 -24626 116 -24593
rect 614 -24626 706 -24593
rect 365 -24626 457 -24593
rect 738 -24626 830 -24593
rect 581 -24626 614 -24593
rect 240 -24626 332 -24593
rect 863 -24626 955 -24593
rect 830 -24768 863 -24735
rect 489 -24768 581 -24735
rect 365 -24768 457 -24735
rect 332 -24768 365 -24735
rect -9 -24768 83 -24735
rect 83 -24768 116 -24735
rect 614 -24768 706 -24735
rect 581 -24768 614 -24735
rect 738 -24768 830 -24735
rect 240 -24768 332 -24735
rect 863 -24768 955 -24735
rect 489 -24910 581 -24877
rect 830 -24910 863 -24877
rect 365 -24910 457 -24877
rect 332 -24910 365 -24877
rect -9 -24910 83 -24877
rect 83 -24910 116 -24877
rect 614 -24910 706 -24877
rect 581 -24910 614 -24877
rect 738 -24910 830 -24877
rect 240 -24910 332 -24877
rect 863 -24910 955 -24877
rect 830 -25052 863 -25019
rect 489 -25052 581 -25019
rect 365 -25052 457 -25019
rect 332 -25052 365 -25019
rect -9 -25052 83 -25019
rect 83 -25052 116 -25019
rect 116 -25052 208 -25019
rect 614 -25052 706 -25019
rect 581 -25052 614 -25019
rect 738 -25052 830 -25019
rect 240 -25052 332 -25019
rect 863 -25052 955 -25019
rect 830 -25194 863 -25161
rect -9 -25194 83 -25161
rect 83 -25194 116 -25161
rect 116 -25194 208 -25161
rect 614 -25194 706 -25161
rect 581 -25194 614 -25161
rect 738 -25194 830 -25161
rect 863 -25194 955 -25161
rect 830 -25336 863 -25303
rect 489 -25336 581 -25303
rect -9 -25336 83 -25303
rect 83 -25336 116 -25303
rect 116 -25336 208 -25303
rect 614 -25336 706 -25303
rect 581 -25336 614 -25303
rect 738 -25336 830 -25303
rect 863 -25336 955 -25303
rect 489 -25478 581 -25445
rect 830 -25478 863 -25445
rect -9 -25478 83 -25445
rect 83 -25478 116 -25445
rect 116 -25478 208 -25445
rect 614 -25478 706 -25445
rect 581 -25478 614 -25445
rect 738 -25478 830 -25445
rect 863 -25478 955 -25445
rect 830 -25620 863 -25587
rect 489 -25620 581 -25587
rect 365 -25620 457 -25587
rect -9 -25620 83 -25587
rect 332 -25620 365 -25587
rect 83 -25620 116 -25587
rect 116 -25620 208 -25587
rect 614 -25620 706 -25587
rect 581 -25620 614 -25587
rect 738 -25620 830 -25587
rect 863 -25620 955 -25587
rect 830 -25762 863 -25729
rect 332 -25762 365 -25729
rect -9 -25762 83 -25729
rect 83 -25762 116 -25729
rect 116 -25762 208 -25729
rect 614 -25762 706 -25729
rect 365 -25762 457 -25729
rect 738 -25762 830 -25729
rect 581 -25762 614 -25729
rect 863 -25762 955 -25729
rect 830 -25904 863 -25871
rect 489 -25904 581 -25871
rect 365 -25904 457 -25871
rect 332 -25904 365 -25871
rect -9 -25904 83 -25871
rect 83 -25904 116 -25871
rect 116 -25904 208 -25871
rect 614 -25904 706 -25871
rect 581 -25904 614 -25871
rect 738 -25904 830 -25871
rect 863 -25904 955 -25871
rect 489 -26046 581 -26013
rect 830 -26046 863 -26013
rect 365 -26046 457 -26013
rect 332 -26046 365 -26013
rect -9 -26046 83 -26013
rect 83 -26046 116 -26013
rect 116 -26046 208 -26013
rect 614 -26046 706 -26013
rect 581 -26046 614 -26013
rect 738 -26046 830 -26013
rect 863 -26046 955 -26013
rect 830 -26188 863 -26155
rect 489 -26188 581 -26155
rect 365 -26188 457 -26155
rect 332 -26188 365 -26155
rect -9 -26188 83 -26155
rect 83 -26188 116 -26155
rect 116 -26188 208 -26155
rect 614 -26188 706 -26155
rect 581 -26188 614 -26155
rect 738 -26188 830 -26155
rect 240 -26188 332 -26155
rect 863 -26188 955 -26155
rect 830 -26330 863 -26297
rect 332 -26330 365 -26297
rect -9 -26330 83 -26297
rect 83 -26330 116 -26297
rect 116 -26330 208 -26297
rect 614 -26330 706 -26297
rect 581 -26330 614 -26297
rect 738 -26330 830 -26297
rect 240 -26330 332 -26297
rect 863 -26330 955 -26297
rect 830 -26472 863 -26439
rect 489 -26472 581 -26439
rect 332 -26472 365 -26439
rect -9 -26472 83 -26439
rect 83 -26472 116 -26439
rect 116 -26472 208 -26439
rect 614 -26472 706 -26439
rect 581 -26472 614 -26439
rect 738 -26472 830 -26439
rect 240 -26472 332 -26439
rect 863 -26472 955 -26439
rect 489 -26614 581 -26581
rect 830 -26614 863 -26581
rect 332 -26614 365 -26581
rect -9 -26614 83 -26581
rect 83 -26614 116 -26581
rect 116 -26614 208 -26581
rect 614 -26614 706 -26581
rect 581 -26614 614 -26581
rect 738 -26614 830 -26581
rect 240 -26614 332 -26581
rect 863 -26614 955 -26581
rect 830 -26756 863 -26723
rect 489 -26756 581 -26723
rect 365 -26756 457 -26723
rect 332 -26756 365 -26723
rect -9 -26756 83 -26723
rect 83 -26756 116 -26723
rect 116 -26756 208 -26723
rect 614 -26756 706 -26723
rect 581 -26756 614 -26723
rect 738 -26756 830 -26723
rect 240 -26756 332 -26723
rect 863 -26756 955 -26723
rect 830 -26898 863 -26865
rect 332 -26898 365 -26865
rect -9 -26898 83 -26865
rect 83 -26898 116 -26865
rect 116 -26898 208 -26865
rect 614 -26898 706 -26865
rect 365 -26898 457 -26865
rect 738 -26898 830 -26865
rect 581 -26898 614 -26865
rect 240 -26898 332 -26865
rect 863 -26898 955 -26865
rect 830 -27040 863 -27007
rect 489 -27040 581 -27007
rect 365 -27040 457 -27007
rect 332 -27040 365 -27007
rect -9 -27040 83 -27007
rect 83 -27040 116 -27007
rect 116 -27040 208 -27007
rect 614 -27040 706 -27007
rect 581 -27040 614 -27007
rect 738 -27040 830 -27007
rect 240 -27040 332 -27007
rect 863 -27040 955 -27007
rect 489 -27182 581 -27149
rect 830 -27182 863 -27149
rect 365 -27182 457 -27149
rect 332 -27182 365 -27149
rect -9 -27182 83 -27149
rect 83 -27182 116 -27149
rect 116 -27182 208 -27149
rect 614 -27182 706 -27149
rect 581 -27182 614 -27149
rect 738 -27182 830 -27149
rect 240 -27182 332 -27149
rect 863 -27182 955 -27149
rect 830 -27324 863 -27291
rect 489 -27324 581 -27291
rect 365 -27324 457 -27291
rect 332 -27324 365 -27291
rect -9 -27324 83 -27291
rect 83 -27324 116 -27291
rect 116 -27324 208 -27291
rect 614 -27324 706 -27291
rect 581 -27324 614 -27291
rect 738 -27324 830 -27291
rect 240 -27324 332 -27291
rect 863 -27324 955 -27291
rect 489 -27466 581 -27433
rect 830 -27466 863 -27433
rect 365 -27466 457 -27433
rect 332 -27466 365 -27433
rect -9 -27466 83 -27433
rect 83 -27466 116 -27433
rect 116 -27466 208 -27433
rect 581 -27466 614 -27433
rect 738 -27466 830 -27433
rect 240 -27466 332 -27433
rect 863 -27466 955 -27433
rect 830 -27608 863 -27575
rect 365 -27608 457 -27575
rect 332 -27608 365 -27575
rect -9 -27608 83 -27575
rect 83 -27608 116 -27575
rect 116 -27608 208 -27575
rect 614 -27608 706 -27575
rect 581 -27608 614 -27575
rect 738 -27608 830 -27575
rect 240 -27608 332 -27575
rect 863 -27608 955 -27575
rect 830 -27750 863 -27717
rect 332 -27750 365 -27717
rect -9 -27750 83 -27717
rect 83 -27750 116 -27717
rect 116 -27750 208 -27717
rect 365 -27750 457 -27717
rect 738 -27750 830 -27717
rect 240 -27750 332 -27717
rect 863 -27750 955 -27717
rect 830 -27892 863 -27859
rect 489 -27892 581 -27859
rect 332 -27892 365 -27859
rect -9 -27892 83 -27859
rect 83 -27892 116 -27859
rect 116 -27892 208 -27859
rect 614 -27892 706 -27859
rect 581 -27892 614 -27859
rect 738 -27892 830 -27859
rect 240 -27892 332 -27859
rect 863 -27892 955 -27859
rect 489 -28034 581 -28001
rect 830 -28034 863 -28001
rect 332 -28034 365 -28001
rect -9 -28034 83 -28001
rect 83 -28034 116 -28001
rect 116 -28034 208 -28001
rect 581 -28034 614 -28001
rect 738 -28034 830 -28001
rect 240 -28034 332 -28001
rect 863 -28034 955 -28001
rect 830 -28176 863 -28143
rect 332 -28176 365 -28143
rect -9 -28176 83 -28143
rect 83 -28176 116 -28143
rect 116 -28176 208 -28143
rect 614 -28176 706 -28143
rect 581 -28176 614 -28143
rect 738 -28176 830 -28143
rect 240 -28176 332 -28143
rect 863 -28176 955 -28143
rect 830 -28318 863 -28285
rect 332 -28318 365 -28285
rect -9 -28318 83 -28285
rect 83 -28318 116 -28285
rect 116 -28318 208 -28285
rect 738 -28318 830 -28285
rect 240 -28318 332 -28285
rect 863 -28318 955 -28285
rect 830 -28460 863 -28427
rect 489 -28460 581 -28427
rect 365 -28460 457 -28427
rect 332 -28460 365 -28427
rect -9 -28460 83 -28427
rect 83 -28460 116 -28427
rect 116 -28460 208 -28427
rect 614 -28460 706 -28427
rect 581 -28460 614 -28427
rect 738 -28460 830 -28427
rect 863 -28460 955 -28427
rect 489 -28602 581 -28569
rect 830 -28602 863 -28569
rect 365 -28602 457 -28569
rect 332 -28602 365 -28569
rect -9 -28602 83 -28569
rect 83 -28602 116 -28569
rect 116 -28602 208 -28569
rect 581 -28602 614 -28569
rect 738 -28602 830 -28569
rect 863 -28602 955 -28569
rect 830 -28744 863 -28711
rect 365 -28744 457 -28711
rect 332 -28744 365 -28711
rect -9 -28744 83 -28711
rect 83 -28744 116 -28711
rect 116 -28744 208 -28711
rect 614 -28744 706 -28711
rect 581 -28744 614 -28711
rect 738 -28744 830 -28711
rect 863 -28744 955 -28711
rect 830 -28886 863 -28853
rect 332 -28886 365 -28853
rect -9 -28886 83 -28853
rect 83 -28886 116 -28853
rect 116 -28886 208 -28853
rect 365 -28886 457 -28853
rect 738 -28886 830 -28853
rect 863 -28886 955 -28853
rect 830 -29028 863 -28995
rect 489 -29028 581 -28995
rect -9 -29028 83 -28995
rect 83 -29028 116 -28995
rect 116 -29028 208 -28995
rect 614 -29028 706 -28995
rect 581 -29028 614 -28995
rect 738 -29028 830 -28995
rect 863 -29028 955 -28995
rect 489 -29170 581 -29137
rect 830 -29170 863 -29137
rect -9 -29170 83 -29137
rect 83 -29170 116 -29137
rect 116 -29170 208 -29137
rect 581 -29170 614 -29137
rect 738 -29170 830 -29137
rect 863 -29170 955 -29137
rect 830 -29312 863 -29279
rect -9 -29312 83 -29279
rect 83 -29312 116 -29279
rect 116 -29312 208 -29279
rect 614 -29312 706 -29279
rect 581 -29312 614 -29279
rect 738 -29312 830 -29279
rect 863 -29312 955 -29279
rect 830 -29454 863 -29421
rect -9 -29454 83 -29421
rect 83 -29454 116 -29421
rect 116 -29454 208 -29421
rect 738 -29454 830 -29421
rect 863 -29454 955 -29421
rect 830 -29596 863 -29563
rect 489 -29596 581 -29563
rect 365 -29596 457 -29563
rect 332 -29596 365 -29563
rect -9 -29596 83 -29563
rect 83 -29596 116 -29563
rect 614 -29596 706 -29563
rect 581 -29596 614 -29563
rect 738 -29596 830 -29563
rect 240 -29596 332 -29563
rect 863 -29596 955 -29563
rect 489 -29738 581 -29705
rect 830 -29738 863 -29705
rect 365 -29738 457 -29705
rect 332 -29738 365 -29705
rect -9 -29738 83 -29705
rect 83 -29738 116 -29705
rect 581 -29738 614 -29705
rect 738 -29738 830 -29705
rect 240 -29738 332 -29705
rect 863 -29738 955 -29705
rect 830 -29880 863 -29847
rect 365 -29880 457 -29847
rect 332 -29880 365 -29847
rect -9 -29880 83 -29847
rect 83 -29880 116 -29847
rect 614 -29880 706 -29847
rect 581 -29880 614 -29847
rect 738 -29880 830 -29847
rect 240 -29880 332 -29847
rect 863 -29880 955 -29847
rect 830 -30022 863 -29989
rect 332 -30022 365 -29989
rect -9 -30022 83 -29989
rect 83 -30022 116 -29989
rect 365 -30022 457 -29989
rect 738 -30022 830 -29989
rect 240 -30022 332 -29989
rect 863 -30022 955 -29989
rect 830 -30164 863 -30131
rect 489 -30164 581 -30131
rect 332 -30164 365 -30131
rect -9 -30164 83 -30131
rect 83 -30164 116 -30131
rect 614 -30164 706 -30131
rect 581 -30164 614 -30131
rect 738 -30164 830 -30131
rect 240 -30164 332 -30131
rect 863 -30164 955 -30131
rect 489 -30306 581 -30273
rect 830 -30306 863 -30273
rect 332 -30306 365 -30273
rect -9 -30306 83 -30273
rect 83 -30306 116 -30273
rect 581 -30306 614 -30273
rect 738 -30306 830 -30273
rect 240 -30306 332 -30273
rect 863 -30306 955 -30273
rect 830 -30448 863 -30415
rect 332 -30448 365 -30415
rect -9 -30448 83 -30415
rect 83 -30448 116 -30415
rect 614 -30448 706 -30415
rect 581 -30448 614 -30415
rect 738 -30448 830 -30415
rect 240 -30448 332 -30415
rect 863 -30448 955 -30415
rect 830 -30590 863 -30557
rect 332 -30590 365 -30557
rect -9 -30590 83 -30557
rect 83 -30590 116 -30557
rect 738 -30590 830 -30557
rect 240 -30590 332 -30557
rect 863 -30590 955 -30557
rect 830 -30732 863 -30699
rect 489 -30732 581 -30699
rect 365 -30732 457 -30699
rect 332 -30732 365 -30699
rect -9 -30732 83 -30699
rect 83 -30732 116 -30699
rect 614 -30732 706 -30699
rect 581 -30732 614 -30699
rect 738 -30732 830 -30699
rect 863 -30732 955 -30699
rect 489 -30874 581 -30841
rect 830 -30874 863 -30841
rect 365 -30874 457 -30841
rect 332 -30874 365 -30841
rect -9 -30874 83 -30841
rect 83 -30874 116 -30841
rect 581 -30874 614 -30841
rect 738 -30874 830 -30841
rect 863 -30874 955 -30841
rect 830 -31016 863 -30983
rect 365 -31016 457 -30983
rect 332 -31016 365 -30983
rect -9 -31016 83 -30983
rect 83 -31016 116 -30983
rect 614 -31016 706 -30983
rect 581 -31016 614 -30983
rect 738 -31016 830 -30983
rect 863 -31016 955 -30983
rect 830 -31158 863 -31125
rect 332 -31158 365 -31125
rect -9 -31158 83 -31125
rect 83 -31158 116 -31125
rect 365 -31158 457 -31125
rect 738 -31158 830 -31125
rect 863 -31158 955 -31125
rect 830 -31300 863 -31267
rect 489 -31300 581 -31267
rect -9 -31300 83 -31267
rect 83 -31300 116 -31267
rect 614 -31300 706 -31267
rect 581 -31300 614 -31267
rect 738 -31300 830 -31267
rect 863 -31300 955 -31267
rect 489 -31442 581 -31409
rect 830 -31442 863 -31409
rect -9 -31442 83 -31409
rect 83 -31442 116 -31409
rect 581 -31442 614 -31409
rect 738 -31442 830 -31409
rect 863 -31442 955 -31409
rect 830 -31584 863 -31551
rect -9 -31584 83 -31551
rect 83 -31584 116 -31551
rect 614 -31584 706 -31551
rect 581 -31584 614 -31551
rect 738 -31584 830 -31551
rect 863 -31584 955 -31551
rect 830 -31726 863 -31693
rect -9 -31726 83 -31693
rect 83 -31726 116 -31693
rect 738 -31726 830 -31693
rect 863 -31726 955 -31693
rect 830 -31868 863 -31835
rect 489 -31868 581 -31835
rect 365 -31868 457 -31835
rect 332 -31868 365 -31835
rect 83 -31868 116 -31835
rect 116 -31868 208 -31835
rect 614 -31868 706 -31835
rect 581 -31868 614 -31835
rect 738 -31868 830 -31835
rect 240 -31868 332 -31835
rect 863 -31868 955 -31835
rect 489 -32010 581 -31977
rect 830 -32010 863 -31977
rect 365 -32010 457 -31977
rect 332 -32010 365 -31977
rect 83 -32010 116 -31977
rect 116 -32010 208 -31977
rect 581 -32010 614 -31977
rect 738 -32010 830 -31977
rect 240 -32010 332 -31977
rect 863 -32010 955 -31977
rect 830 -32152 863 -32119
rect 365 -32152 457 -32119
rect 332 -32152 365 -32119
rect 83 -32152 116 -32119
rect 116 -32152 208 -32119
rect 614 -32152 706 -32119
rect 581 -32152 614 -32119
rect 738 -32152 830 -32119
rect 240 -32152 332 -32119
rect 863 -32152 955 -32119
rect 830 -32294 863 -32261
rect 332 -32294 365 -32261
rect 83 -32294 116 -32261
rect 116 -32294 208 -32261
rect 365 -32294 457 -32261
rect 738 -32294 830 -32261
rect 240 -32294 332 -32261
rect 863 -32294 955 -32261
rect 830 -32436 863 -32403
rect 489 -32436 581 -32403
rect 332 -32436 365 -32403
rect 83 -32436 116 -32403
rect 116 -32436 208 -32403
rect 614 -32436 706 -32403
rect 581 -32436 614 -32403
rect 738 -32436 830 -32403
rect 240 -32436 332 -32403
rect 863 -32436 955 -32403
rect 489 -32578 581 -32545
rect 830 -32578 863 -32545
rect 332 -32578 365 -32545
rect 83 -32578 116 -32545
rect 116 -32578 208 -32545
rect 581 -32578 614 -32545
rect 738 -32578 830 -32545
rect 240 -32578 332 -32545
rect 863 -32578 955 -32545
rect 830 -32720 863 -32687
rect 332 -32720 365 -32687
rect 83 -32720 116 -32687
rect 116 -32720 208 -32687
rect 614 -32720 706 -32687
rect 581 -32720 614 -32687
rect 738 -32720 830 -32687
rect 240 -32720 332 -32687
rect 863 -32720 955 -32687
rect 830 -32862 863 -32829
rect 332 -32862 365 -32829
rect 83 -32862 116 -32829
rect 116 -32862 208 -32829
rect 738 -32862 830 -32829
rect 240 -32862 332 -32829
rect 863 -32862 955 -32829
rect 830 -33004 863 -32971
rect 489 -33004 581 -32971
rect 365 -33004 457 -32971
rect 332 -33004 365 -32971
rect 83 -33004 116 -32971
rect 116 -33004 208 -32971
rect 614 -33004 706 -32971
rect 581 -33004 614 -32971
rect 738 -33004 830 -32971
rect 863 -33004 955 -32971
rect 489 -33146 581 -33113
rect 830 -33146 863 -33113
rect 365 -33146 457 -33113
rect 332 -33146 365 -33113
rect 83 -33146 116 -33113
rect 116 -33146 208 -33113
rect 581 -33146 614 -33113
rect 738 -33146 830 -33113
rect 863 -33146 955 -33113
rect 830 -33288 863 -33255
rect 365 -33288 457 -33255
rect 332 -33288 365 -33255
rect 83 -33288 116 -33255
rect 116 -33288 208 -33255
rect 614 -33288 706 -33255
rect 581 -33288 614 -33255
rect 738 -33288 830 -33255
rect 863 -33288 955 -33255
rect 830 -33430 863 -33397
rect 332 -33430 365 -33397
rect 83 -33430 116 -33397
rect 116 -33430 208 -33397
rect 365 -33430 457 -33397
rect 738 -33430 830 -33397
rect 863 -33430 955 -33397
rect 830 -33572 863 -33539
rect 489 -33572 581 -33539
rect 83 -33572 116 -33539
rect 116 -33572 208 -33539
rect 614 -33572 706 -33539
rect 581 -33572 614 -33539
rect 738 -33572 830 -33539
rect 863 -33572 955 -33539
rect 489 -33714 581 -33681
rect 830 -33714 863 -33681
rect 83 -33714 116 -33681
rect 116 -33714 208 -33681
rect 581 -33714 614 -33681
rect 738 -33714 830 -33681
rect 863 -33714 955 -33681
rect 830 -33856 863 -33823
rect 83 -33856 116 -33823
rect 116 -33856 208 -33823
rect 614 -33856 706 -33823
rect 581 -33856 614 -33823
rect 738 -33856 830 -33823
rect 863 -33856 955 -33823
rect 830 -33998 863 -33965
rect 83 -33998 116 -33965
rect 116 -33998 208 -33965
rect 738 -33998 830 -33965
rect 863 -33998 955 -33965
rect 830 -34140 863 -34107
rect 489 -34140 581 -34107
rect 365 -34140 457 -34107
rect 332 -34140 365 -34107
rect 614 -34140 706 -34107
rect 581 -34140 614 -34107
rect 738 -34140 830 -34107
rect 240 -34140 332 -34107
rect 863 -34140 955 -34107
rect 489 -34282 581 -34249
rect 830 -34282 863 -34249
rect 365 -34282 457 -34249
rect 332 -34282 365 -34249
rect 581 -34282 614 -34249
rect 738 -34282 830 -34249
rect 240 -34282 332 -34249
rect 863 -34282 955 -34249
rect 830 -34424 863 -34391
rect 365 -34424 457 -34391
rect 332 -34424 365 -34391
rect 614 -34424 706 -34391
rect 581 -34424 614 -34391
rect 738 -34424 830 -34391
rect 240 -34424 332 -34391
rect 863 -34424 955 -34391
rect 830 -34566 863 -34533
rect 332 -34566 365 -34533
rect 365 -34566 457 -34533
rect 738 -34566 830 -34533
rect 240 -34566 332 -34533
rect 863 -34566 955 -34533
rect 830 -34708 863 -34675
rect 489 -34708 581 -34675
rect 332 -34708 365 -34675
rect 614 -34708 706 -34675
rect 581 -34708 614 -34675
rect 738 -34708 830 -34675
rect 240 -34708 332 -34675
rect 863 -34708 955 -34675
rect 489 -34850 581 -34817
rect 830 -34850 863 -34817
rect 332 -34850 365 -34817
rect 581 -34850 614 -34817
rect 738 -34850 830 -34817
rect 240 -34850 332 -34817
rect 863 -34850 955 -34817
rect 830 -34992 863 -34959
rect 332 -34992 365 -34959
rect 614 -34992 706 -34959
rect 581 -34992 614 -34959
rect 738 -34992 830 -34959
rect 240 -34992 332 -34959
rect 863 -34992 955 -34959
rect 830 -35134 863 -35101
rect 332 -35134 365 -35101
rect 738 -35134 830 -35101
rect 240 -35134 332 -35101
rect 863 -35134 955 -35101
rect 830 -35276 863 -35243
rect 489 -35276 581 -35243
rect 365 -35276 457 -35243
rect 332 -35276 365 -35243
rect 614 -35276 706 -35243
rect 581 -35276 614 -35243
rect 738 -35276 830 -35243
rect 863 -35276 955 -35243
rect 489 -35418 581 -35385
rect 830 -35418 863 -35385
rect 365 -35418 457 -35385
rect 332 -35418 365 -35385
rect 581 -35418 614 -35385
rect 738 -35418 830 -35385
rect 863 -35418 955 -35385
rect 830 -35560 863 -35527
rect 365 -35560 457 -35527
rect 332 -35560 365 -35527
rect 614 -35560 706 -35527
rect 581 -35560 614 -35527
rect 738 -35560 830 -35527
rect 863 -35560 955 -35527
rect 830 -35702 863 -35669
rect 332 -35702 365 -35669
rect 365 -35702 457 -35669
rect 738 -35702 830 -35669
rect 863 -35702 955 -35669
rect 830 -35844 863 -35811
rect 489 -35844 581 -35811
rect 614 -35844 706 -35811
rect 581 -35844 614 -35811
rect 738 -35844 830 -35811
rect 863 -35844 955 -35811
rect 489 -35986 581 -35953
rect 830 -35986 863 -35953
rect 581 -35986 614 -35953
rect 738 -35986 830 -35953
rect 863 -35986 955 -35953
rect 830 -36128 863 -36095
rect 614 -36128 706 -36095
rect 581 -36128 614 -36095
rect 738 -36128 830 -36095
rect 863 -36128 955 -36095
rect 738 -36270 830 -36237
rect 830 -36270 863 -36237
rect 863 -36270 955 -36237
rect 738 -36554 830 -36521
rect 830 -36554 863 -36521
rect 863 -36554 955 -36521
rect 830 -36696 863 -36663
rect 614 -36696 706 -36663
rect 581 -36696 614 -36663
rect 738 -36696 830 -36663
rect 863 -36696 955 -36663
rect 830 -36838 863 -36805
rect 614 -36838 706 -36805
rect 581 -36838 614 -36805
rect 738 -36838 830 -36805
rect 863 -36838 955 -36805
rect 830 -36980 863 -36947
rect 489 -36980 581 -36947
rect 614 -36980 706 -36947
rect 581 -36980 614 -36947
rect 738 -36980 830 -36947
rect 863 -36980 955 -36947
rect 489 -37122 581 -37089
rect 830 -37122 863 -37089
rect 581 -37122 614 -37089
rect 738 -37122 830 -37089
rect 863 -37122 955 -37089
rect 489 -37264 581 -37231
rect 830 -37264 863 -37231
rect 614 -37264 706 -37231
rect 581 -37264 614 -37231
rect 738 -37264 830 -37231
rect 863 -37264 955 -37231
rect 489 -37406 581 -37373
rect 830 -37406 863 -37373
rect 614 -37406 706 -37373
rect 581 -37406 614 -37373
rect 738 -37406 830 -37373
rect 863 -37406 955 -37373
rect 830 -37548 863 -37515
rect 489 -37548 581 -37515
rect 365 -37548 457 -37515
rect 332 -37548 365 -37515
rect 614 -37548 706 -37515
rect 581 -37548 614 -37515
rect 738 -37548 830 -37515
rect 863 -37548 955 -37515
rect 830 -37690 863 -37657
rect 332 -37690 365 -37657
rect 365 -37690 457 -37657
rect 738 -37690 830 -37657
rect 863 -37690 955 -37657
rect 830 -37832 863 -37799
rect 332 -37832 365 -37799
rect 614 -37832 706 -37799
rect 365 -37832 457 -37799
rect 738 -37832 830 -37799
rect 581 -37832 614 -37799
rect 863 -37832 955 -37799
rect 830 -37974 863 -37941
rect 365 -37974 457 -37941
rect 332 -37974 365 -37941
rect 614 -37974 706 -37941
rect 581 -37974 614 -37941
rect 738 -37974 830 -37941
rect 863 -37974 955 -37941
rect 830 -38116 863 -38083
rect 489 -38116 581 -38083
rect 365 -38116 457 -38083
rect 332 -38116 365 -38083
rect 614 -38116 706 -38083
rect 581 -38116 614 -38083
rect 738 -38116 830 -38083
rect 863 -38116 955 -38083
rect 489 -38258 581 -38225
rect 830 -38258 863 -38225
rect 365 -38258 457 -38225
rect 332 -38258 365 -38225
rect 581 -38258 614 -38225
rect 738 -38258 830 -38225
rect 863 -38258 955 -38225
rect 489 -38400 581 -38367
rect 830 -38400 863 -38367
rect 365 -38400 457 -38367
rect 332 -38400 365 -38367
rect 614 -38400 706 -38367
rect 581 -38400 614 -38367
rect 738 -38400 830 -38367
rect 863 -38400 955 -38367
rect 489 -38542 581 -38509
rect 830 -38542 863 -38509
rect 365 -38542 457 -38509
rect 332 -38542 365 -38509
rect 614 -38542 706 -38509
rect 581 -38542 614 -38509
rect 738 -38542 830 -38509
rect 863 -38542 955 -38509
rect 830 -38684 863 -38651
rect 489 -38684 581 -38651
rect 365 -38684 457 -38651
rect 332 -38684 365 -38651
rect 614 -38684 706 -38651
rect 581 -38684 614 -38651
rect 738 -38684 830 -38651
rect 240 -38684 332 -38651
rect 863 -38684 955 -38651
rect 830 -38826 863 -38793
rect 332 -38826 365 -38793
rect 738 -38826 830 -38793
rect 240 -38826 332 -38793
rect 863 -38826 955 -38793
rect 830 -38968 863 -38935
rect 332 -38968 365 -38935
rect 614 -38968 706 -38935
rect 581 -38968 614 -38935
rect 738 -38968 830 -38935
rect 240 -38968 332 -38935
rect 863 -38968 955 -38935
rect 830 -39110 863 -39077
rect 332 -39110 365 -39077
rect 614 -39110 706 -39077
rect 581 -39110 614 -39077
rect 738 -39110 830 -39077
rect 240 -39110 332 -39077
rect 863 -39110 955 -39077
rect 830 -39252 863 -39219
rect 489 -39252 581 -39219
rect 332 -39252 365 -39219
rect 614 -39252 706 -39219
rect 581 -39252 614 -39219
rect 738 -39252 830 -39219
rect 240 -39252 332 -39219
rect 863 -39252 955 -39219
rect 489 -39394 581 -39361
rect 830 -39394 863 -39361
rect 332 -39394 365 -39361
rect 581 -39394 614 -39361
rect 738 -39394 830 -39361
rect 240 -39394 332 -39361
rect 863 -39394 955 -39361
rect 489 -39536 581 -39503
rect 830 -39536 863 -39503
rect 332 -39536 365 -39503
rect 614 -39536 706 -39503
rect 581 -39536 614 -39503
rect 738 -39536 830 -39503
rect 240 -39536 332 -39503
rect 863 -39536 955 -39503
rect 489 -39678 581 -39645
rect 830 -39678 863 -39645
rect 332 -39678 365 -39645
rect 614 -39678 706 -39645
rect 581 -39678 614 -39645
rect 738 -39678 830 -39645
rect 240 -39678 332 -39645
rect 863 -39678 955 -39645
rect 830 -39820 863 -39787
rect 489 -39820 581 -39787
rect 365 -39820 457 -39787
rect 332 -39820 365 -39787
rect 614 -39820 706 -39787
rect 581 -39820 614 -39787
rect 738 -39820 830 -39787
rect 240 -39820 332 -39787
rect 863 -39820 955 -39787
rect 830 -39962 863 -39929
rect 332 -39962 365 -39929
rect 365 -39962 457 -39929
rect 738 -39962 830 -39929
rect 240 -39962 332 -39929
rect 863 -39962 955 -39929
rect 830 -40104 863 -40071
rect 332 -40104 365 -40071
rect 614 -40104 706 -40071
rect 365 -40104 457 -40071
rect 738 -40104 830 -40071
rect 581 -40104 614 -40071
rect 240 -40104 332 -40071
rect 863 -40104 955 -40071
rect 830 -40246 863 -40213
rect 365 -40246 457 -40213
rect 332 -40246 365 -40213
rect 614 -40246 706 -40213
rect 581 -40246 614 -40213
rect 738 -40246 830 -40213
rect 240 -40246 332 -40213
rect 863 -40246 955 -40213
rect 830 -40388 863 -40355
rect 489 -40388 581 -40355
rect 365 -40388 457 -40355
rect 332 -40388 365 -40355
rect 614 -40388 706 -40355
rect 581 -40388 614 -40355
rect 738 -40388 830 -40355
rect 240 -40388 332 -40355
rect 863 -40388 955 -40355
rect 489 -40530 581 -40497
rect 830 -40530 863 -40497
rect 365 -40530 457 -40497
rect 332 -40530 365 -40497
rect 581 -40530 614 -40497
rect 738 -40530 830 -40497
rect 240 -40530 332 -40497
rect 863 -40530 955 -40497
rect 489 -40672 581 -40639
rect 830 -40672 863 -40639
rect 365 -40672 457 -40639
rect 332 -40672 365 -40639
rect 614 -40672 706 -40639
rect 581 -40672 614 -40639
rect 738 -40672 830 -40639
rect 240 -40672 332 -40639
rect 863 -40672 955 -40639
rect 489 -40814 581 -40781
rect 830 -40814 863 -40781
rect 365 -40814 457 -40781
rect 332 -40814 365 -40781
rect 614 -40814 706 -40781
rect 581 -40814 614 -40781
rect 738 -40814 830 -40781
rect 240 -40814 332 -40781
rect 863 -40814 955 -40781
rect 830 -40956 863 -40923
rect 489 -40956 581 -40923
rect 365 -40956 457 -40923
rect 332 -40956 365 -40923
rect 83 -40956 116 -40923
rect 116 -40956 208 -40923
rect 614 -40956 706 -40923
rect 581 -40956 614 -40923
rect 738 -40956 830 -40923
rect 240 -40956 332 -40923
rect 863 -40956 955 -40923
rect 830 -41098 863 -41065
rect 83 -41098 116 -41065
rect 116 -41098 208 -41065
rect 738 -41098 830 -41065
rect 863 -41098 955 -41065
rect 830 -41240 863 -41207
rect 83 -41240 116 -41207
rect 116 -41240 208 -41207
rect 614 -41240 706 -41207
rect 581 -41240 614 -41207
rect 738 -41240 830 -41207
rect 863 -41240 955 -41207
rect 830 -41382 863 -41349
rect 83 -41382 116 -41349
rect 116 -41382 208 -41349
rect 614 -41382 706 -41349
rect 581 -41382 614 -41349
rect 738 -41382 830 -41349
rect 863 -41382 955 -41349
rect 830 -41524 863 -41491
rect 489 -41524 581 -41491
rect 83 -41524 116 -41491
rect 116 -41524 208 -41491
rect 614 -41524 706 -41491
rect 581 -41524 614 -41491
rect 738 -41524 830 -41491
rect 863 -41524 955 -41491
rect 489 -41666 581 -41633
rect 830 -41666 863 -41633
rect 83 -41666 116 -41633
rect 116 -41666 208 -41633
rect 581 -41666 614 -41633
rect 738 -41666 830 -41633
rect 863 -41666 955 -41633
rect 489 -41808 581 -41775
rect 830 -41808 863 -41775
rect 83 -41808 116 -41775
rect 116 -41808 208 -41775
rect 614 -41808 706 -41775
rect 581 -41808 614 -41775
rect 738 -41808 830 -41775
rect 863 -41808 955 -41775
rect 489 -41950 581 -41917
rect 830 -41950 863 -41917
rect 83 -41950 116 -41917
rect 116 -41950 208 -41917
rect 614 -41950 706 -41917
rect 581 -41950 614 -41917
rect 738 -41950 830 -41917
rect 863 -41950 955 -41917
rect 830 -42092 863 -42059
rect 489 -42092 581 -42059
rect 365 -42092 457 -42059
rect 332 -42092 365 -42059
rect 83 -42092 116 -42059
rect 116 -42092 208 -42059
rect 614 -42092 706 -42059
rect 581 -42092 614 -42059
rect 738 -42092 830 -42059
rect 863 -42092 955 -42059
rect 830 -42234 863 -42201
rect 332 -42234 365 -42201
rect 83 -42234 116 -42201
rect 116 -42234 208 -42201
rect 365 -42234 457 -42201
rect 738 -42234 830 -42201
rect 863 -42234 955 -42201
rect 830 -42376 863 -42343
rect 332 -42376 365 -42343
rect 83 -42376 116 -42343
rect 116 -42376 208 -42343
rect 614 -42376 706 -42343
rect 365 -42376 457 -42343
rect 738 -42376 830 -42343
rect 581 -42376 614 -42343
rect 863 -42376 955 -42343
rect 830 -42518 863 -42485
rect 365 -42518 457 -42485
rect 332 -42518 365 -42485
rect 83 -42518 116 -42485
rect 116 -42518 208 -42485
rect 614 -42518 706 -42485
rect 581 -42518 614 -42485
rect 738 -42518 830 -42485
rect 863 -42518 955 -42485
rect 830 -42660 863 -42627
rect 489 -42660 581 -42627
rect 365 -42660 457 -42627
rect 332 -42660 365 -42627
rect 83 -42660 116 -42627
rect 116 -42660 208 -42627
rect 614 -42660 706 -42627
rect 581 -42660 614 -42627
rect 738 -42660 830 -42627
rect 863 -42660 955 -42627
rect 489 -42802 581 -42769
rect 830 -42802 863 -42769
rect 365 -42802 457 -42769
rect 332 -42802 365 -42769
rect 83 -42802 116 -42769
rect 116 -42802 208 -42769
rect 581 -42802 614 -42769
rect 738 -42802 830 -42769
rect 863 -42802 955 -42769
rect 489 -42944 581 -42911
rect 830 -42944 863 -42911
rect 365 -42944 457 -42911
rect 332 -42944 365 -42911
rect 83 -42944 116 -42911
rect 116 -42944 208 -42911
rect 614 -42944 706 -42911
rect 581 -42944 614 -42911
rect 738 -42944 830 -42911
rect 863 -42944 955 -42911
rect 489 -43086 581 -43053
rect 830 -43086 863 -43053
rect 365 -43086 457 -43053
rect 332 -43086 365 -43053
rect 83 -43086 116 -43053
rect 116 -43086 208 -43053
rect 614 -43086 706 -43053
rect 581 -43086 614 -43053
rect 738 -43086 830 -43053
rect 863 -43086 955 -43053
rect 830 -43228 863 -43195
rect 489 -43228 581 -43195
rect 365 -43228 457 -43195
rect 332 -43228 365 -43195
rect 83 -43228 116 -43195
rect 116 -43228 208 -43195
rect 614 -43228 706 -43195
rect 581 -43228 614 -43195
rect 738 -43228 830 -43195
rect 240 -43228 332 -43195
rect 863 -43228 955 -43195
rect 830 -43370 863 -43337
rect 332 -43370 365 -43337
rect 83 -43370 116 -43337
rect 116 -43370 208 -43337
rect 738 -43370 830 -43337
rect 240 -43370 332 -43337
rect 863 -43370 955 -43337
rect 830 -43512 863 -43479
rect 332 -43512 365 -43479
rect 83 -43512 116 -43479
rect 116 -43512 208 -43479
rect 614 -43512 706 -43479
rect 581 -43512 614 -43479
rect 738 -43512 830 -43479
rect 240 -43512 332 -43479
rect 863 -43512 955 -43479
rect 830 -43654 863 -43621
rect 332 -43654 365 -43621
rect 83 -43654 116 -43621
rect 116 -43654 208 -43621
rect 614 -43654 706 -43621
rect 581 -43654 614 -43621
rect 738 -43654 830 -43621
rect 240 -43654 332 -43621
rect 863 -43654 955 -43621
rect 830 -43796 863 -43763
rect 489 -43796 581 -43763
rect 332 -43796 365 -43763
rect 83 -43796 116 -43763
rect 116 -43796 208 -43763
rect 614 -43796 706 -43763
rect 581 -43796 614 -43763
rect 738 -43796 830 -43763
rect 240 -43796 332 -43763
rect 863 -43796 955 -43763
rect 489 -43938 581 -43905
rect 830 -43938 863 -43905
rect 332 -43938 365 -43905
rect 83 -43938 116 -43905
rect 116 -43938 208 -43905
rect 581 -43938 614 -43905
rect 738 -43938 830 -43905
rect 240 -43938 332 -43905
rect 863 -43938 955 -43905
rect 489 -44080 581 -44047
rect 830 -44080 863 -44047
rect 332 -44080 365 -44047
rect 83 -44080 116 -44047
rect 116 -44080 208 -44047
rect 614 -44080 706 -44047
rect 581 -44080 614 -44047
rect 738 -44080 830 -44047
rect 240 -44080 332 -44047
rect 863 -44080 955 -44047
rect 489 -44222 581 -44189
rect 830 -44222 863 -44189
rect 332 -44222 365 -44189
rect 83 -44222 116 -44189
rect 116 -44222 208 -44189
rect 614 -44222 706 -44189
rect 581 -44222 614 -44189
rect 738 -44222 830 -44189
rect 240 -44222 332 -44189
rect 863 -44222 955 -44189
rect 830 -44364 863 -44331
rect 489 -44364 581 -44331
rect 365 -44364 457 -44331
rect 332 -44364 365 -44331
rect 83 -44364 116 -44331
rect 116 -44364 208 -44331
rect 614 -44364 706 -44331
rect 581 -44364 614 -44331
rect 738 -44364 830 -44331
rect 240 -44364 332 -44331
rect 863 -44364 955 -44331
rect 830 -44506 863 -44473
rect 332 -44506 365 -44473
rect 83 -44506 116 -44473
rect 116 -44506 208 -44473
rect 365 -44506 457 -44473
rect 738 -44506 830 -44473
rect 240 -44506 332 -44473
rect 863 -44506 955 -44473
rect 830 -44648 863 -44615
rect 332 -44648 365 -44615
rect 83 -44648 116 -44615
rect 116 -44648 208 -44615
rect 614 -44648 706 -44615
rect 365 -44648 457 -44615
rect 738 -44648 830 -44615
rect 581 -44648 614 -44615
rect 240 -44648 332 -44615
rect 863 -44648 955 -44615
rect 830 -44790 863 -44757
rect 365 -44790 457 -44757
rect 332 -44790 365 -44757
rect 83 -44790 116 -44757
rect 116 -44790 208 -44757
rect 614 -44790 706 -44757
rect 581 -44790 614 -44757
rect 738 -44790 830 -44757
rect 240 -44790 332 -44757
rect 863 -44790 955 -44757
rect 830 -44932 863 -44899
rect 489 -44932 581 -44899
rect 365 -44932 457 -44899
rect 332 -44932 365 -44899
rect 83 -44932 116 -44899
rect 116 -44932 208 -44899
rect 614 -44932 706 -44899
rect 581 -44932 614 -44899
rect 738 -44932 830 -44899
rect 240 -44932 332 -44899
rect 863 -44932 955 -44899
rect 489 -45074 581 -45041
rect 830 -45074 863 -45041
rect 365 -45074 457 -45041
rect 332 -45074 365 -45041
rect 83 -45074 116 -45041
rect 116 -45074 208 -45041
rect 581 -45074 614 -45041
rect 738 -45074 830 -45041
rect 240 -45074 332 -45041
rect 863 -45074 955 -45041
rect 489 -45216 581 -45183
rect 830 -45216 863 -45183
rect 365 -45216 457 -45183
rect 332 -45216 365 -45183
rect 83 -45216 116 -45183
rect 116 -45216 208 -45183
rect 614 -45216 706 -45183
rect 581 -45216 614 -45183
rect 738 -45216 830 -45183
rect 240 -45216 332 -45183
rect 863 -45216 955 -45183
rect 489 -45358 581 -45325
rect 830 -45358 863 -45325
rect 365 -45358 457 -45325
rect 332 -45358 365 -45325
rect 83 -45358 116 -45325
rect 116 -45358 208 -45325
rect 614 -45358 706 -45325
rect 581 -45358 614 -45325
rect 738 -45358 830 -45325
rect 240 -45358 332 -45325
rect 863 -45358 955 -45325
rect 830 -45500 863 -45467
rect 489 -45500 581 -45467
rect 365 -45500 457 -45467
rect 332 -45500 365 -45467
rect -9 -45500 83 -45467
rect 83 -45500 116 -45467
rect 116 -45500 208 -45467
rect 614 -45500 706 -45467
rect 581 -45500 614 -45467
rect 738 -45500 830 -45467
rect 240 -45500 332 -45467
rect 863 -45500 955 -45467
rect 830 -45642 863 -45609
rect -9 -45642 83 -45609
rect 83 -45642 116 -45609
rect 738 -45642 830 -45609
rect 863 -45642 955 -45609
rect 830 -45784 863 -45751
rect -9 -45784 83 -45751
rect 83 -45784 116 -45751
rect 614 -45784 706 -45751
rect 581 -45784 614 -45751
rect 738 -45784 830 -45751
rect 863 -45784 955 -45751
rect 830 -45926 863 -45893
rect -9 -45926 83 -45893
rect 83 -45926 116 -45893
rect 614 -45926 706 -45893
rect 581 -45926 614 -45893
rect 738 -45926 830 -45893
rect 863 -45926 955 -45893
rect 830 -46068 863 -46035
rect 489 -46068 581 -46035
rect -9 -46068 83 -46035
rect 83 -46068 116 -46035
rect 614 -46068 706 -46035
rect 581 -46068 614 -46035
rect 738 -46068 830 -46035
rect 863 -46068 955 -46035
rect 489 -46210 581 -46177
rect 830 -46210 863 -46177
rect -9 -46210 83 -46177
rect 83 -46210 116 -46177
rect 581 -46210 614 -46177
rect 738 -46210 830 -46177
rect 863 -46210 955 -46177
rect 489 -46352 581 -46319
rect 830 -46352 863 -46319
rect -9 -46352 83 -46319
rect 83 -46352 116 -46319
rect 614 -46352 706 -46319
rect 581 -46352 614 -46319
rect 738 -46352 830 -46319
rect 863 -46352 955 -46319
rect 489 -46494 581 -46461
rect 830 -46494 863 -46461
rect -9 -46494 83 -46461
rect 83 -46494 116 -46461
rect 614 -46494 706 -46461
rect 581 -46494 614 -46461
rect 738 -46494 830 -46461
rect 863 -46494 955 -46461
rect 830 -46636 863 -46603
rect 489 -46636 581 -46603
rect 365 -46636 457 -46603
rect -9 -46636 83 -46603
rect 332 -46636 365 -46603
rect 83 -46636 116 -46603
rect 614 -46636 706 -46603
rect 581 -46636 614 -46603
rect 738 -46636 830 -46603
rect 863 -46636 955 -46603
rect 830 -46778 863 -46745
rect 332 -46778 365 -46745
rect -9 -46778 83 -46745
rect 83 -46778 116 -46745
rect 365 -46778 457 -46745
rect 738 -46778 830 -46745
rect 863 -46778 955 -46745
rect 830 -46920 863 -46887
rect 332 -46920 365 -46887
rect -9 -46920 83 -46887
rect 83 -46920 116 -46887
rect 614 -46920 706 -46887
rect 365 -46920 457 -46887
rect 738 -46920 830 -46887
rect 581 -46920 614 -46887
rect 863 -46920 955 -46887
rect 830 -47062 863 -47029
rect 365 -47062 457 -47029
rect 332 -47062 365 -47029
rect -9 -47062 83 -47029
rect 83 -47062 116 -47029
rect 614 -47062 706 -47029
rect 581 -47062 614 -47029
rect 738 -47062 830 -47029
rect 863 -47062 955 -47029
rect 830 -47204 863 -47171
rect 489 -47204 581 -47171
rect 365 -47204 457 -47171
rect 332 -47204 365 -47171
rect -9 -47204 83 -47171
rect 83 -47204 116 -47171
rect 614 -47204 706 -47171
rect 581 -47204 614 -47171
rect 738 -47204 830 -47171
rect 863 -47204 955 -47171
rect 489 -47346 581 -47313
rect 830 -47346 863 -47313
rect 365 -47346 457 -47313
rect 332 -47346 365 -47313
rect -9 -47346 83 -47313
rect 83 -47346 116 -47313
rect 581 -47346 614 -47313
rect 738 -47346 830 -47313
rect 863 -47346 955 -47313
rect 489 -47488 581 -47455
rect 830 -47488 863 -47455
rect 365 -47488 457 -47455
rect 332 -47488 365 -47455
rect -9 -47488 83 -47455
rect 83 -47488 116 -47455
rect 614 -47488 706 -47455
rect 581 -47488 614 -47455
rect 738 -47488 830 -47455
rect 863 -47488 955 -47455
rect 489 -47630 581 -47597
rect 830 -47630 863 -47597
rect 365 -47630 457 -47597
rect 332 -47630 365 -47597
rect -9 -47630 83 -47597
rect 83 -47630 116 -47597
rect 614 -47630 706 -47597
rect 581 -47630 614 -47597
rect 738 -47630 830 -47597
rect 863 -47630 955 -47597
rect 830 -47772 863 -47739
rect 489 -47772 581 -47739
rect 365 -47772 457 -47739
rect 332 -47772 365 -47739
rect -9 -47772 83 -47739
rect 83 -47772 116 -47739
rect 614 -47772 706 -47739
rect 581 -47772 614 -47739
rect 738 -47772 830 -47739
rect 240 -47772 332 -47739
rect 863 -47772 955 -47739
rect 830 -47914 863 -47881
rect 332 -47914 365 -47881
rect -9 -47914 83 -47881
rect 83 -47914 116 -47881
rect 738 -47914 830 -47881
rect 240 -47914 332 -47881
rect 863 -47914 955 -47881
rect 830 -48056 863 -48023
rect 332 -48056 365 -48023
rect -9 -48056 83 -48023
rect 83 -48056 116 -48023
rect 614 -48056 706 -48023
rect 581 -48056 614 -48023
rect 738 -48056 830 -48023
rect 240 -48056 332 -48023
rect 863 -48056 955 -48023
rect 830 -48198 863 -48165
rect 332 -48198 365 -48165
rect -9 -48198 83 -48165
rect 83 -48198 116 -48165
rect 614 -48198 706 -48165
rect 581 -48198 614 -48165
rect 738 -48198 830 -48165
rect 240 -48198 332 -48165
rect 863 -48198 955 -48165
rect 830 -48340 863 -48307
rect 489 -48340 581 -48307
rect 332 -48340 365 -48307
rect -9 -48340 83 -48307
rect 83 -48340 116 -48307
rect 614 -48340 706 -48307
rect 581 -48340 614 -48307
rect 738 -48340 830 -48307
rect 240 -48340 332 -48307
rect 863 -48340 955 -48307
rect 489 -48482 581 -48449
rect 830 -48482 863 -48449
rect 332 -48482 365 -48449
rect -9 -48482 83 -48449
rect 83 -48482 116 -48449
rect 581 -48482 614 -48449
rect 738 -48482 830 -48449
rect 240 -48482 332 -48449
rect 863 -48482 955 -48449
rect 489 -48624 581 -48591
rect 830 -48624 863 -48591
rect 332 -48624 365 -48591
rect -9 -48624 83 -48591
rect 83 -48624 116 -48591
rect 614 -48624 706 -48591
rect 581 -48624 614 -48591
rect 738 -48624 830 -48591
rect 240 -48624 332 -48591
rect 863 -48624 955 -48591
rect 489 -48766 581 -48733
rect 830 -48766 863 -48733
rect 332 -48766 365 -48733
rect -9 -48766 83 -48733
rect 83 -48766 116 -48733
rect 614 -48766 706 -48733
rect 581 -48766 614 -48733
rect 738 -48766 830 -48733
rect 240 -48766 332 -48733
rect 863 -48766 955 -48733
rect 830 -48908 863 -48875
rect 489 -48908 581 -48875
rect 365 -48908 457 -48875
rect 332 -48908 365 -48875
rect -9 -48908 83 -48875
rect 83 -48908 116 -48875
rect 614 -48908 706 -48875
rect 581 -48908 614 -48875
rect 738 -48908 830 -48875
rect 240 -48908 332 -48875
rect 863 -48908 955 -48875
rect 830 -49050 863 -49017
rect 332 -49050 365 -49017
rect -9 -49050 83 -49017
rect 83 -49050 116 -49017
rect 365 -49050 457 -49017
rect 738 -49050 830 -49017
rect 240 -49050 332 -49017
rect 863 -49050 955 -49017
rect 830 -49192 863 -49159
rect 332 -49192 365 -49159
rect -9 -49192 83 -49159
rect 83 -49192 116 -49159
rect 614 -49192 706 -49159
rect 365 -49192 457 -49159
rect 738 -49192 830 -49159
rect 581 -49192 614 -49159
rect 240 -49192 332 -49159
rect 863 -49192 955 -49159
rect 830 -49334 863 -49301
rect 365 -49334 457 -49301
rect 332 -49334 365 -49301
rect -9 -49334 83 -49301
rect 83 -49334 116 -49301
rect 614 -49334 706 -49301
rect 581 -49334 614 -49301
rect 738 -49334 830 -49301
rect 240 -49334 332 -49301
rect 863 -49334 955 -49301
rect 830 -49476 863 -49443
rect 489 -49476 581 -49443
rect 365 -49476 457 -49443
rect 332 -49476 365 -49443
rect -9 -49476 83 -49443
rect 83 -49476 116 -49443
rect 614 -49476 706 -49443
rect 581 -49476 614 -49443
rect 738 -49476 830 -49443
rect 240 -49476 332 -49443
rect 863 -49476 955 -49443
rect 489 -49618 581 -49585
rect 830 -49618 863 -49585
rect 365 -49618 457 -49585
rect 332 -49618 365 -49585
rect -9 -49618 83 -49585
rect 83 -49618 116 -49585
rect 581 -49618 614 -49585
rect 738 -49618 830 -49585
rect 240 -49618 332 -49585
rect 863 -49618 955 -49585
rect 489 -49760 581 -49727
rect 830 -49760 863 -49727
rect 365 -49760 457 -49727
rect 332 -49760 365 -49727
rect -9 -49760 83 -49727
rect 83 -49760 116 -49727
rect 614 -49760 706 -49727
rect 581 -49760 614 -49727
rect 738 -49760 830 -49727
rect 240 -49760 332 -49727
rect 863 -49760 955 -49727
rect 489 -49902 581 -49869
rect 830 -49902 863 -49869
rect 365 -49902 457 -49869
rect 332 -49902 365 -49869
rect -9 -49902 83 -49869
rect 83 -49902 116 -49869
rect 614 -49902 706 -49869
rect 581 -49902 614 -49869
rect 738 -49902 830 -49869
rect 240 -49902 332 -49869
rect 863 -49902 955 -49869
rect 830 -50044 863 -50011
rect 489 -50044 581 -50011
rect 365 -50044 457 -50011
rect 332 -50044 365 -50011
rect -9 -50044 83 -50011
rect 83 -50044 116 -50011
rect 116 -50044 208 -50011
rect 614 -50044 706 -50011
rect 581 -50044 614 -50011
rect 738 -50044 830 -50011
rect 240 -50044 332 -50011
rect 863 -50044 955 -50011
rect 830 -50186 863 -50153
rect -9 -50186 83 -50153
rect 83 -50186 116 -50153
rect 116 -50186 208 -50153
rect 738 -50186 830 -50153
rect 863 -50186 955 -50153
rect 830 -50328 863 -50295
rect -9 -50328 83 -50295
rect 83 -50328 116 -50295
rect 116 -50328 208 -50295
rect 614 -50328 706 -50295
rect 581 -50328 614 -50295
rect 738 -50328 830 -50295
rect 863 -50328 955 -50295
rect 830 -50470 863 -50437
rect -9 -50470 83 -50437
rect 83 -50470 116 -50437
rect 116 -50470 208 -50437
rect 614 -50470 706 -50437
rect 581 -50470 614 -50437
rect 738 -50470 830 -50437
rect 863 -50470 955 -50437
rect 830 -50612 863 -50579
rect 489 -50612 581 -50579
rect -9 -50612 83 -50579
rect 83 -50612 116 -50579
rect 116 -50612 208 -50579
rect 614 -50612 706 -50579
rect 581 -50612 614 -50579
rect 738 -50612 830 -50579
rect 863 -50612 955 -50579
rect 489 -50754 581 -50721
rect 830 -50754 863 -50721
rect -9 -50754 83 -50721
rect 83 -50754 116 -50721
rect 116 -50754 208 -50721
rect 581 -50754 614 -50721
rect 738 -50754 830 -50721
rect 863 -50754 955 -50721
rect 489 -50896 581 -50863
rect 830 -50896 863 -50863
rect -9 -50896 83 -50863
rect 83 -50896 116 -50863
rect 116 -50896 208 -50863
rect 614 -50896 706 -50863
rect 581 -50896 614 -50863
rect 738 -50896 830 -50863
rect 863 -50896 955 -50863
rect 489 -51038 581 -51005
rect 830 -51038 863 -51005
rect -9 -51038 83 -51005
rect 83 -51038 116 -51005
rect 116 -51038 208 -51005
rect 614 -51038 706 -51005
rect 581 -51038 614 -51005
rect 738 -51038 830 -51005
rect 863 -51038 955 -51005
rect 830 -51180 863 -51147
rect 489 -51180 581 -51147
rect 365 -51180 457 -51147
rect -9 -51180 83 -51147
rect 332 -51180 365 -51147
rect 83 -51180 116 -51147
rect 116 -51180 208 -51147
rect 614 -51180 706 -51147
rect 581 -51180 614 -51147
rect 738 -51180 830 -51147
rect 863 -51180 955 -51147
rect 830 -51322 863 -51289
rect 332 -51322 365 -51289
rect -9 -51322 83 -51289
rect 83 -51322 116 -51289
rect 116 -51322 208 -51289
rect 365 -51322 457 -51289
rect 738 -51322 830 -51289
rect 863 -51322 955 -51289
rect 830 -51464 863 -51431
rect 332 -51464 365 -51431
rect -9 -51464 83 -51431
rect 83 -51464 116 -51431
rect 116 -51464 208 -51431
rect 614 -51464 706 -51431
rect 365 -51464 457 -51431
rect 738 -51464 830 -51431
rect 581 -51464 614 -51431
rect 863 -51464 955 -51431
rect 830 -51606 863 -51573
rect 365 -51606 457 -51573
rect 332 -51606 365 -51573
rect -9 -51606 83 -51573
rect 83 -51606 116 -51573
rect 116 -51606 208 -51573
rect 614 -51606 706 -51573
rect 581 -51606 614 -51573
rect 738 -51606 830 -51573
rect 863 -51606 955 -51573
rect 830 -51748 863 -51715
rect 489 -51748 581 -51715
rect 365 -51748 457 -51715
rect 332 -51748 365 -51715
rect -9 -51748 83 -51715
rect 83 -51748 116 -51715
rect 116 -51748 208 -51715
rect 614 -51748 706 -51715
rect 581 -51748 614 -51715
rect 738 -51748 830 -51715
rect 863 -51748 955 -51715
rect 489 -51890 581 -51857
rect 830 -51890 863 -51857
rect 365 -51890 457 -51857
rect 332 -51890 365 -51857
rect -9 -51890 83 -51857
rect 83 -51890 116 -51857
rect 116 -51890 208 -51857
rect 581 -51890 614 -51857
rect 738 -51890 830 -51857
rect 863 -51890 955 -51857
rect 489 -52032 581 -51999
rect 830 -52032 863 -51999
rect 365 -52032 457 -51999
rect 332 -52032 365 -51999
rect -9 -52032 83 -51999
rect 83 -52032 116 -51999
rect 116 -52032 208 -51999
rect 614 -52032 706 -51999
rect 581 -52032 614 -51999
rect 738 -52032 830 -51999
rect 863 -52032 955 -51999
rect 489 -52174 581 -52141
rect 830 -52174 863 -52141
rect 365 -52174 457 -52141
rect 332 -52174 365 -52141
rect -9 -52174 83 -52141
rect 83 -52174 116 -52141
rect 116 -52174 208 -52141
rect 614 -52174 706 -52141
rect 581 -52174 614 -52141
rect 738 -52174 830 -52141
rect 863 -52174 955 -52141
rect 830 -52316 863 -52283
rect 489 -52316 581 -52283
rect 365 -52316 457 -52283
rect 332 -52316 365 -52283
rect -9 -52316 83 -52283
rect 83 -52316 116 -52283
rect 116 -52316 208 -52283
rect 614 -52316 706 -52283
rect 581 -52316 614 -52283
rect 738 -52316 830 -52283
rect 240 -52316 332 -52283
rect 863 -52316 955 -52283
rect 830 -52458 863 -52425
rect 332 -52458 365 -52425
rect -9 -52458 83 -52425
rect 83 -52458 116 -52425
rect 116 -52458 208 -52425
rect 738 -52458 830 -52425
rect 240 -52458 332 -52425
rect 863 -52458 955 -52425
rect 830 -52600 863 -52567
rect 332 -52600 365 -52567
rect -9 -52600 83 -52567
rect 83 -52600 116 -52567
rect 116 -52600 208 -52567
rect 614 -52600 706 -52567
rect 581 -52600 614 -52567
rect 738 -52600 830 -52567
rect 240 -52600 332 -52567
rect 863 -52600 955 -52567
rect 830 -52742 863 -52709
rect 332 -52742 365 -52709
rect -9 -52742 83 -52709
rect 83 -52742 116 -52709
rect 116 -52742 208 -52709
rect 614 -52742 706 -52709
rect 581 -52742 614 -52709
rect 738 -52742 830 -52709
rect 240 -52742 332 -52709
rect 863 -52742 955 -52709
rect 830 -52884 863 -52851
rect 489 -52884 581 -52851
rect 332 -52884 365 -52851
rect -9 -52884 83 -52851
rect 83 -52884 116 -52851
rect 116 -52884 208 -52851
rect 614 -52884 706 -52851
rect 581 -52884 614 -52851
rect 738 -52884 830 -52851
rect 240 -52884 332 -52851
rect 863 -52884 955 -52851
rect 489 -53026 581 -52993
rect 830 -53026 863 -52993
rect 332 -53026 365 -52993
rect -9 -53026 83 -52993
rect 83 -53026 116 -52993
rect 116 -53026 208 -52993
rect 581 -53026 614 -52993
rect 738 -53026 830 -52993
rect 240 -53026 332 -52993
rect 863 -53026 955 -52993
rect 489 -53168 581 -53135
rect 830 -53168 863 -53135
rect 332 -53168 365 -53135
rect -9 -53168 83 -53135
rect 83 -53168 116 -53135
rect 116 -53168 208 -53135
rect 614 -53168 706 -53135
rect 581 -53168 614 -53135
rect 738 -53168 830 -53135
rect 240 -53168 332 -53135
rect 863 -53168 955 -53135
rect 489 -53310 581 -53277
rect 830 -53310 863 -53277
rect 332 -53310 365 -53277
rect -9 -53310 83 -53277
rect 83 -53310 116 -53277
rect 116 -53310 208 -53277
rect 614 -53310 706 -53277
rect 581 -53310 614 -53277
rect 738 -53310 830 -53277
rect 240 -53310 332 -53277
rect 863 -53310 955 -53277
rect 830 -53452 863 -53419
rect 489 -53452 581 -53419
rect 365 -53452 457 -53419
rect 332 -53452 365 -53419
rect -9 -53452 83 -53419
rect 83 -53452 116 -53419
rect 116 -53452 208 -53419
rect 614 -53452 706 -53419
rect 581 -53452 614 -53419
rect 738 -53452 830 -53419
rect 240 -53452 332 -53419
rect 863 -53452 955 -53419
rect 830 -53594 863 -53561
rect 332 -53594 365 -53561
rect -9 -53594 83 -53561
rect 83 -53594 116 -53561
rect 116 -53594 208 -53561
rect 365 -53594 457 -53561
rect 738 -53594 830 -53561
rect 240 -53594 332 -53561
rect 863 -53594 955 -53561
rect 830 -53736 863 -53703
rect 332 -53736 365 -53703
rect -9 -53736 83 -53703
rect 83 -53736 116 -53703
rect 116 -53736 208 -53703
rect 614 -53736 706 -53703
rect 365 -53736 457 -53703
rect 738 -53736 830 -53703
rect 581 -53736 614 -53703
rect 240 -53736 332 -53703
rect 863 -53736 955 -53703
rect 830 -53878 863 -53845
rect 365 -53878 457 -53845
rect 332 -53878 365 -53845
rect -9 -53878 83 -53845
rect 83 -53878 116 -53845
rect 116 -53878 208 -53845
rect 614 -53878 706 -53845
rect 581 -53878 614 -53845
rect 738 -53878 830 -53845
rect 240 -53878 332 -53845
rect 863 -53878 955 -53845
rect 830 -54020 863 -53987
rect 489 -54020 581 -53987
rect 365 -54020 457 -53987
rect 332 -54020 365 -53987
rect -9 -54020 83 -53987
rect 83 -54020 116 -53987
rect 116 -54020 208 -53987
rect 614 -54020 706 -53987
rect 581 -54020 614 -53987
rect 738 -54020 830 -53987
rect 240 -54020 332 -53987
rect 863 -54020 955 -53987
rect 489 -54162 581 -54129
rect 830 -54162 863 -54129
rect 365 -54162 457 -54129
rect 332 -54162 365 -54129
rect -9 -54162 83 -54129
rect 83 -54162 116 -54129
rect 116 -54162 208 -54129
rect 581 -54162 614 -54129
rect 738 -54162 830 -54129
rect 240 -54162 332 -54129
rect 863 -54162 955 -54129
rect 489 -54304 581 -54271
rect 830 -54304 863 -54271
rect 365 -54304 457 -54271
rect 332 -54304 365 -54271
rect -9 -54304 83 -54271
rect 83 -54304 116 -54271
rect 116 -54304 208 -54271
rect 614 -54304 706 -54271
rect 581 -54304 614 -54271
rect 738 -54304 830 -54271
rect 240 -54304 332 -54271
rect 863 -54304 955 -54271
rect 489 -54446 581 -54413
rect 830 -54446 863 -54413
rect 365 -54446 457 -54413
rect 332 -54446 365 -54413
rect -9 -54446 83 -54413
rect 83 -54446 116 -54413
rect 116 -54446 208 -54413
rect 614 -54446 706 -54413
rect 581 -54446 614 -54413
rect 738 -54446 830 -54413
rect 240 -54446 332 -54413
rect 863 -54446 955 -54413
rect 830 -54872 863 -54839
rect 863 -54872 955 -54839
rect 738 -55014 830 -54981
rect 830 -55014 863 -54981
rect 863 -55014 955 -54981
rect 738 -55156 830 -55123
rect 830 -55156 863 -55123
rect 863 -55156 955 -55123
rect 581 -55298 614 -55265
rect 863 -55298 955 -55265
rect 830 -55298 863 -55265
rect 614 -55298 706 -55265
rect 830 -55440 863 -55407
rect 614 -55440 706 -55407
rect 581 -55440 614 -55407
rect 738 -55440 830 -55407
rect 863 -55440 955 -55407
rect 830 -55582 863 -55549
rect 489 -55582 581 -55549
rect 614 -55582 706 -55549
rect 581 -55582 614 -55549
rect 738 -55582 830 -55549
rect 863 -55582 955 -55549
rect 489 -55724 581 -55691
rect 830 -55724 863 -55691
rect 581 -55724 614 -55691
rect 738 -55724 830 -55691
rect 863 -55724 955 -55691
rect 830 -55866 863 -55833
rect 489 -55866 581 -55833
rect 614 -55866 706 -55833
rect 581 -55866 614 -55833
rect 738 -55866 830 -55833
rect 830 -56008 863 -55975
rect 489 -56008 581 -55975
rect 365 -56008 457 -55975
rect 332 -56008 365 -55975
rect 614 -56008 706 -55975
rect 581 -56008 614 -55975
rect 738 -56008 830 -55975
rect 863 -56008 955 -55975
rect 830 -56150 863 -56117
rect 332 -56150 365 -56117
rect 614 -56150 706 -56117
rect 365 -56150 457 -56117
rect 738 -56150 830 -56117
rect 581 -56150 614 -56117
rect 830 -56292 863 -56259
rect 365 -56292 457 -56259
rect 332 -56292 365 -56259
rect 614 -56292 706 -56259
rect 581 -56292 614 -56259
rect 738 -56292 830 -56259
rect 863 -56292 955 -56259
rect 489 -56434 581 -56401
rect 830 -56434 863 -56401
rect 365 -56434 457 -56401
rect 332 -56434 365 -56401
rect 581 -56434 614 -56401
rect 738 -56434 830 -56401
rect 863 -56434 955 -56401
rect 489 -56576 581 -56543
rect 830 -56576 863 -56543
rect 365 -56576 457 -56543
rect 332 -56576 365 -56543
rect 614 -56576 706 -56543
rect 581 -56576 614 -56543
rect 738 -56576 830 -56543
rect 863 -56576 955 -56543
rect 830 -56718 863 -56685
rect 332 -56718 365 -56685
rect 738 -56718 830 -56685
rect 240 -56718 332 -56685
rect 863 -56718 955 -56685
rect 830 -56860 863 -56827
rect 489 -56860 581 -56827
rect 332 -56860 365 -56827
rect 614 -56860 706 -56827
rect 581 -56860 614 -56827
rect 240 -56860 332 -56827
rect 863 -56860 955 -56827
rect 489 -57002 581 -56969
rect 830 -57002 863 -56969
rect 332 -57002 365 -56969
rect 614 -57002 706 -56969
rect 581 -57002 614 -56969
rect 738 -57002 830 -56969
rect 240 -57002 332 -56969
rect 830 -57144 863 -57111
rect 489 -57144 581 -57111
rect 365 -57144 457 -57111
rect 332 -57144 365 -57111
rect 614 -57144 706 -57111
rect 581 -57144 614 -57111
rect 738 -57144 830 -57111
rect 240 -57144 332 -57111
rect 863 -57144 955 -57111
rect 830 -57286 863 -57253
rect 365 -57286 457 -57253
rect 332 -57286 365 -57253
rect 614 -57286 706 -57253
rect 581 -57286 614 -57253
rect 738 -57286 830 -57253
rect 240 -57286 332 -57253
rect 489 -57428 581 -57395
rect 830 -57428 863 -57395
rect 365 -57428 457 -57395
rect 332 -57428 365 -57395
rect 581 -57428 614 -57395
rect 738 -57428 830 -57395
rect 240 -57428 332 -57395
rect 863 -57428 955 -57395
rect 489 -57570 581 -57537
rect 830 -57570 863 -57537
rect 365 -57570 457 -57537
rect 332 -57570 365 -57537
rect 83 -57570 116 -57537
rect 116 -57570 208 -57537
rect 614 -57570 706 -57537
rect 581 -57570 614 -57537
rect 738 -57570 830 -57537
rect 240 -57570 332 -57537
rect 863 -57570 955 -57537
rect 830 -57712 863 -57679
rect 83 -57712 116 -57679
rect 116 -57712 208 -57679
rect 614 -57712 706 -57679
rect 581 -57712 614 -57679
rect 738 -57712 830 -57679
rect 863 -57712 955 -57679
rect 489 -57854 581 -57821
rect 830 -57854 863 -57821
rect 83 -57854 116 -57821
rect 116 -57854 208 -57821
rect 614 -57854 706 -57821
rect 581 -57854 614 -57821
rect 863 -57854 955 -57821
rect 830 -57996 863 -57963
rect 489 -57996 581 -57963
rect 365 -57996 457 -57963
rect 332 -57996 365 -57963
rect 83 -57996 116 -57963
rect 116 -57996 208 -57963
rect 614 -57996 706 -57963
rect 581 -57996 614 -57963
rect 738 -57996 830 -57963
rect 863 -57996 955 -57963
rect 830 -58138 863 -58105
rect 489 -58138 581 -58105
rect 365 -58138 457 -58105
rect 332 -58138 365 -58105
rect 83 -58138 116 -58105
rect 116 -58138 208 -58105
rect 614 -58138 706 -58105
rect 581 -58138 614 -58105
rect 863 -58138 955 -58105
rect 489 -58280 581 -58247
rect 830 -58280 863 -58247
rect 365 -58280 457 -58247
rect 332 -58280 365 -58247
rect 83 -58280 116 -58247
rect 116 -58280 208 -58247
rect 614 -58280 706 -58247
rect 581 -58280 614 -58247
rect 738 -58280 830 -58247
rect 863 -58280 955 -58247
rect 830 -58422 863 -58389
rect 332 -58422 365 -58389
rect 83 -58422 116 -58389
rect 116 -58422 208 -58389
rect 614 -58422 706 -58389
rect 581 -58422 614 -58389
rect 240 -58422 332 -58389
rect 863 -58422 955 -58389
rect 830 -58564 863 -58531
rect 489 -58564 581 -58531
rect 332 -58564 365 -58531
rect 83 -58564 116 -58531
rect 116 -58564 208 -58531
rect 614 -58564 706 -58531
rect 581 -58564 614 -58531
rect 738 -58564 830 -58531
rect 240 -58564 332 -58531
rect 863 -58564 955 -58531
rect 489 -58706 581 -58673
rect 830 -58706 863 -58673
rect 365 -58706 457 -58673
rect 332 -58706 365 -58673
rect 83 -58706 116 -58673
rect 116 -58706 208 -58673
rect 614 -58706 706 -58673
rect 581 -58706 614 -58673
rect 240 -58706 332 -58673
rect 863 -58706 955 -58673
rect 830 -58848 863 -58815
rect 332 -58848 365 -58815
rect 83 -58848 116 -58815
rect 116 -58848 208 -58815
rect 614 -58848 706 -58815
rect 365 -58848 457 -58815
rect 738 -58848 830 -58815
rect 581 -58848 614 -58815
rect 240 -58848 332 -58815
rect 863 -58848 955 -58815
rect 489 -58990 581 -58957
rect 830 -58990 863 -58957
rect 365 -58990 457 -58957
rect 332 -58990 365 -58957
rect 83 -58990 116 -58957
rect 116 -58990 208 -58957
rect 614 -58990 706 -58957
rect 581 -58990 614 -58957
rect 240 -58990 332 -58957
rect 863 -58990 955 -58957
rect 830 -59132 863 -59099
rect -9 -59132 83 -59099
rect 83 -59132 116 -59099
rect 738 -59132 830 -59099
rect 863 -59132 955 -59099
rect 830 -59274 863 -59241
rect 489 -59274 581 -59241
rect -9 -59274 83 -59241
rect 83 -59274 116 -59241
rect 614 -59274 706 -59241
rect 581 -59274 614 -59241
rect 738 -59274 830 -59241
rect 863 -59274 955 -59241
rect 489 -59416 581 -59383
rect 830 -59416 863 -59383
rect -9 -59416 83 -59383
rect 83 -59416 116 -59383
rect 614 -59416 706 -59383
rect 581 -59416 614 -59383
rect 738 -59416 830 -59383
rect 863 -59416 955 -59383
rect 830 -59558 863 -59525
rect 332 -59558 365 -59525
rect -9 -59558 83 -59525
rect 83 -59558 116 -59525
rect 614 -59558 706 -59525
rect 365 -59558 457 -59525
rect 738 -59558 830 -59525
rect 581 -59558 614 -59525
rect 863 -59558 955 -59525
rect 489 -59700 581 -59667
rect 830 -59700 863 -59667
rect 365 -59700 457 -59667
rect 332 -59700 365 -59667
rect -9 -59700 83 -59667
rect 83 -59700 116 -59667
rect 581 -59700 614 -59667
rect 738 -59700 830 -59667
rect 863 -59700 955 -59667
rect 489 -59842 581 -59809
rect 830 -59842 863 -59809
rect 365 -59842 457 -59809
rect 332 -59842 365 -59809
rect -9 -59842 83 -59809
rect 83 -59842 116 -59809
rect 614 -59842 706 -59809
rect 581 -59842 614 -59809
rect 738 -59842 830 -59809
rect 240 -59842 332 -59809
rect 830 -59984 863 -59951
rect 332 -59984 365 -59951
rect -9 -59984 83 -59951
rect 83 -59984 116 -59951
rect 614 -59984 706 -59951
rect 581 -59984 614 -59951
rect 738 -59984 830 -59951
rect 240 -59984 332 -59951
rect 863 -59984 955 -59951
rect 489 -60126 581 -60093
rect 830 -60126 863 -60093
rect 332 -60126 365 -60093
rect -9 -60126 83 -60093
rect 83 -60126 116 -60093
rect 614 -60126 706 -60093
rect 581 -60126 614 -60093
rect 738 -60126 830 -60093
rect 240 -60126 332 -60093
rect 863 -60126 955 -60093
rect 830 -60268 863 -60235
rect 332 -60268 365 -60235
rect -9 -60268 83 -60235
rect 83 -60268 116 -60235
rect 365 -60268 457 -60235
rect 738 -60268 830 -60235
rect 240 -60268 332 -60235
rect 863 -60268 955 -60235
rect 830 -60410 863 -60377
rect 489 -60410 581 -60377
rect 365 -60410 457 -60377
rect 332 -60410 365 -60377
rect -9 -60410 83 -60377
rect 83 -60410 116 -60377
rect 614 -60410 706 -60377
rect 581 -60410 614 -60377
rect 738 -60410 830 -60377
rect 240 -60410 332 -60377
rect 863 -60410 955 -60377
rect 489 -60552 581 -60519
rect 830 -60552 863 -60519
rect 365 -60552 457 -60519
rect 332 -60552 365 -60519
rect -9 -60552 83 -60519
rect 83 -60552 116 -60519
rect 614 -60552 706 -60519
rect 581 -60552 614 -60519
rect 738 -60552 830 -60519
rect 240 -60552 332 -60519
rect 830 -60694 863 -60661
rect -9 -60694 83 -60661
rect 83 -60694 116 -60661
rect 116 -60694 208 -60661
rect 614 -60694 706 -60661
rect 581 -60694 614 -60661
rect 863 -60694 955 -60661
rect 830 -60836 863 -60803
rect 489 -60836 581 -60803
rect -9 -60836 83 -60803
rect 83 -60836 116 -60803
rect 116 -60836 208 -60803
rect 614 -60836 706 -60803
rect 581 -60836 614 -60803
rect 738 -60836 830 -60803
rect 863 -60836 955 -60803
rect 489 -60978 581 -60945
rect 830 -60978 863 -60945
rect -9 -60978 83 -60945
rect 83 -60978 116 -60945
rect 116 -60978 208 -60945
rect 614 -60978 706 -60945
rect 581 -60978 614 -60945
rect 738 -60978 830 -60945
rect 863 -60978 955 -60945
rect 830 -61120 863 -61087
rect 332 -61120 365 -61087
rect -9 -61120 83 -61087
rect 83 -61120 116 -61087
rect 116 -61120 208 -61087
rect 365 -61120 457 -61087
rect 738 -61120 830 -61087
rect 863 -61120 955 -61087
rect 830 -61262 863 -61229
rect 365 -61262 457 -61229
rect 332 -61262 365 -61229
rect -9 -61262 83 -61229
rect 83 -61262 116 -61229
rect 116 -61262 208 -61229
rect 614 -61262 706 -61229
rect 581 -61262 614 -61229
rect 738 -61262 830 -61229
rect 863 -61262 955 -61229
rect 489 -61404 581 -61371
rect 830 -61404 863 -61371
rect 365 -61404 457 -61371
rect 332 -61404 365 -61371
rect -9 -61404 83 -61371
rect 83 -61404 116 -61371
rect 116 -61404 208 -61371
rect 614 -61404 706 -61371
rect 581 -61404 614 -61371
rect 738 -61404 830 -61371
rect 489 -61546 581 -61513
rect 830 -61546 863 -61513
rect 365 -61546 457 -61513
rect 332 -61546 365 -61513
rect -9 -61546 83 -61513
rect 83 -61546 116 -61513
rect 116 -61546 208 -61513
rect 614 -61546 706 -61513
rect 581 -61546 614 -61513
rect 738 -61546 830 -61513
rect 240 -61546 332 -61513
rect 830 -61688 863 -61655
rect 332 -61688 365 -61655
rect -9 -61688 83 -61655
rect 83 -61688 116 -61655
rect 116 -61688 208 -61655
rect 614 -61688 706 -61655
rect 581 -61688 614 -61655
rect 738 -61688 830 -61655
rect 240 -61688 332 -61655
rect 830 -61830 863 -61797
rect 489 -61830 581 -61797
rect 332 -61830 365 -61797
rect -9 -61830 83 -61797
rect 83 -61830 116 -61797
rect 116 -61830 208 -61797
rect 614 -61830 706 -61797
rect 581 -61830 614 -61797
rect 738 -61830 830 -61797
rect 240 -61830 332 -61797
rect 489 -61972 581 -61939
rect 830 -61972 863 -61939
rect 332 -61972 365 -61939
rect -9 -61972 83 -61939
rect 83 -61972 116 -61939
rect 116 -61972 208 -61939
rect 581 -61972 614 -61939
rect 738 -61972 830 -61939
rect 240 -61972 332 -61939
rect 863 -61972 955 -61939
rect 489 -62114 581 -62081
rect 830 -62114 863 -62081
rect 332 -62114 365 -62081
rect -9 -62114 83 -62081
rect 83 -62114 116 -62081
rect 116 -62114 208 -62081
rect 614 -62114 706 -62081
rect 581 -62114 614 -62081
rect 738 -62114 830 -62081
rect 240 -62114 332 -62081
rect 863 -62114 955 -62081
rect 830 -62256 863 -62223
rect 332 -62256 365 -62223
rect -9 -62256 83 -62223
rect 83 -62256 116 -62223
rect 116 -62256 208 -62223
rect 365 -62256 457 -62223
rect 240 -62256 332 -62223
rect 863 -62256 955 -62223
rect 830 -62398 863 -62365
rect 332 -62398 365 -62365
rect -9 -62398 83 -62365
rect 83 -62398 116 -62365
rect 116 -62398 208 -62365
rect 614 -62398 706 -62365
rect 365 -62398 457 -62365
rect 738 -62398 830 -62365
rect 581 -62398 614 -62365
rect 240 -62398 332 -62365
rect 863 -62398 955 -62365
rect 830 -62540 863 -62507
rect 365 -62540 457 -62507
rect 332 -62540 365 -62507
rect -9 -62540 83 -62507
rect 83 -62540 116 -62507
rect 116 -62540 208 -62507
rect 614 -62540 706 -62507
rect 581 -62540 614 -62507
rect 738 -62540 830 -62507
rect 240 -62540 332 -62507
rect 863 -62540 955 -62507
rect 489 -62682 581 -62649
rect 830 -62682 863 -62649
rect 365 -62682 457 -62649
rect 332 -62682 365 -62649
rect -9 -62682 83 -62649
rect 83 -62682 116 -62649
rect 116 -62682 208 -62649
rect 581 -62682 614 -62649
rect 240 -62682 332 -62649
rect 863 -62682 955 -62649
rect 489 -62824 581 -62791
rect 830 -62824 863 -62791
rect 365 -62824 457 -62791
rect 332 -62824 365 -62791
rect -9 -62824 83 -62791
rect 83 -62824 116 -62791
rect 116 -62824 208 -62791
rect 581 -62824 614 -62791
rect 738 -62824 830 -62791
rect 240 -62824 332 -62791
rect 489 -62966 581 -62933
rect 830 -62966 863 -62933
rect 365 -62966 457 -62933
rect 332 -62966 365 -62933
rect -9 -62966 83 -62933
rect 83 -62966 116 -62933
rect 116 -62966 208 -62933
rect 614 -62966 706 -62933
rect 581 -62966 614 -62933
rect 738 -62966 830 -62933
rect 240 -62966 332 -62933
rect 863 -62966 955 -62933
rect 489 -63108 581 -63075
rect 830 -63108 863 -63075
rect 365 -63108 457 -63075
rect 332 -63108 365 -63075
rect -9 -63108 83 -63075
rect 83 -63108 116 -63075
rect 116 -63108 208 -63075
rect 614 -63108 706 -63075
rect 581 -63108 614 -63075
rect 240 -63108 332 -63075
rect 863 -63108 955 -63075
rect 489 -63250 581 -63217
rect 830 -63250 863 -63217
rect 365 -63250 457 -63217
rect 332 -63250 365 -63217
rect -9 -63250 83 -63217
rect 83 -63250 116 -63217
rect 116 -63250 208 -63217
rect 614 -63250 706 -63217
rect 581 -63250 614 -63217
rect 738 -63250 830 -63217
rect 240 -63250 332 -63217
rect 489 -63392 581 -63359
rect 830 -63392 863 -63359
rect 365 -63392 457 -63359
rect 332 -63392 365 -63359
rect -9 -63392 83 -63359
rect 83 -63392 116 -63359
rect 116 -63392 208 -63359
rect 614 -63392 706 -63359
rect 581 -63392 614 -63359
rect 738 -63392 830 -63359
rect 240 -63392 332 -63359
rect 863 -63392 955 -63359
rect 830 -63534 863 -63501
rect 489 -63534 581 -63501
rect 365 -63534 457 -63501
rect 332 -63534 365 -63501
rect -9 -63534 83 -63501
rect 83 -63534 116 -63501
rect 116 -63534 208 -63501
rect 614 -63534 706 -63501
rect 581 -63534 614 -63501
rect 738 -63534 830 -63501
rect 240 -63534 332 -63501
rect 863 -63534 955 -63501
rect 830 -63676 863 -63643
rect 489 -63676 581 -63643
rect 365 -63676 457 -63643
rect 332 -63676 365 -63643
rect -9 -63676 83 -63643
rect 83 -63676 116 -63643
rect 116 -63676 208 -63643
rect 614 -63676 706 -63643
rect 581 -63676 614 -63643
rect 738 -63676 830 -63643
rect 240 -63676 332 -63643
rect 863 -63676 955 -63643
rect 830 -63818 863 -63785
rect 489 -63818 581 -63785
rect 365 -63818 457 -63785
rect 332 -63818 365 -63785
rect -9 -63818 83 -63785
rect 83 -63818 116 -63785
rect 116 -63818 208 -63785
rect 614 -63818 706 -63785
rect 581 -63818 614 -63785
rect 738 -63818 830 -63785
rect 240 -63818 332 -63785
rect 863 -63818 955 -63785
rect 489 -63960 581 -63927
rect 830 -63960 863 -63927
rect 365 -63960 457 -63927
rect 332 -63960 365 -63927
rect -9 -63960 83 -63927
rect 83 -63960 116 -63927
rect 116 -63960 208 -63927
rect 614 -63960 706 -63927
rect 581 -63960 614 -63927
rect 738 -63960 830 -63927
rect 240 -63960 332 -63927
rect 489 -64102 581 -64069
rect 830 -64102 863 -64069
rect 365 -64102 457 -64069
rect 332 -64102 365 -64069
rect -9 -64102 83 -64069
rect 83 -64102 116 -64069
rect 116 -64102 208 -64069
rect 614 -64102 706 -64069
rect 581 -64102 614 -64069
rect 738 -64102 830 -64069
rect 240 -64102 332 -64069
rect 863 -64102 955 -64069
rect 489 -64244 581 -64211
rect 830 -64244 863 -64211
rect 365 -64244 457 -64211
rect 332 -64244 365 -64211
rect -9 -64244 83 -64211
rect 83 -64244 116 -64211
rect 116 -64244 208 -64211
rect 614 -64244 706 -64211
rect 581 -64244 614 -64211
rect 240 -64244 332 -64211
rect 863 -64244 955 -64211
rect 489 -64386 581 -64353
rect 830 -64386 863 -64353
rect 365 -64386 457 -64353
rect 332 -64386 365 -64353
rect -9 -64386 83 -64353
rect 83 -64386 116 -64353
rect 116 -64386 208 -64353
rect 581 -64386 614 -64353
rect 738 -64386 830 -64353
rect 240 -64386 332 -64353
rect 863 -64386 955 -64353
rect 489 -64528 581 -64495
rect 830 -64528 863 -64495
rect 365 -64528 457 -64495
rect 332 -64528 365 -64495
rect -9 -64528 83 -64495
rect 83 -64528 116 -64495
rect 116 -64528 208 -64495
rect 581 -64528 614 -64495
rect 738 -64528 830 -64495
rect 240 -64528 332 -64495
rect 863 -64528 955 -64495
rect 489 -64670 581 -64637
rect 830 -64670 863 -64637
rect 365 -64670 457 -64637
rect 332 -64670 365 -64637
rect -9 -64670 83 -64637
rect 83 -64670 116 -64637
rect 116 -64670 208 -64637
rect 614 -64670 706 -64637
rect 581 -64670 614 -64637
rect 738 -64670 830 -64637
rect 240 -64670 332 -64637
rect 830 -64812 863 -64779
rect 365 -64812 457 -64779
rect 332 -64812 365 -64779
rect -9 -64812 83 -64779
rect 83 -64812 116 -64779
rect 116 -64812 208 -64779
rect 614 -64812 706 -64779
rect 581 -64812 614 -64779
rect 240 -64812 332 -64779
rect 863 -64812 955 -64779
rect 830 -64954 863 -64921
rect 332 -64954 365 -64921
rect -9 -64954 83 -64921
rect 83 -64954 116 -64921
rect 116 -64954 208 -64921
rect 365 -64954 457 -64921
rect 738 -64954 830 -64921
rect 240 -64954 332 -64921
rect 863 -64954 955 -64921
rect 830 -65096 863 -65063
rect 489 -65096 581 -65063
rect 332 -65096 365 -65063
rect -9 -65096 83 -65063
rect 83 -65096 116 -65063
rect 116 -65096 208 -65063
rect 614 -65096 706 -65063
rect 365 -65096 457 -65063
rect 738 -65096 830 -65063
rect 581 -65096 614 -65063
rect 240 -65096 332 -65063
rect 489 -65238 581 -65205
rect 830 -65238 863 -65205
rect 332 -65238 365 -65205
rect -9 -65238 83 -65205
rect 83 -65238 116 -65205
rect 116 -65238 208 -65205
rect 614 -65238 706 -65205
rect 581 -65238 614 -65205
rect 738 -65238 830 -65205
rect 240 -65238 332 -65205
rect 863 -65238 955 -65205
rect 489 -65380 581 -65347
rect 830 -65380 863 -65347
rect 332 -65380 365 -65347
rect -9 -65380 83 -65347
rect 83 -65380 116 -65347
rect 116 -65380 208 -65347
rect 581 -65380 614 -65347
rect 738 -65380 830 -65347
rect 240 -65380 332 -65347
rect 830 -65522 863 -65489
rect 332 -65522 365 -65489
rect -9 -65522 83 -65489
rect 83 -65522 116 -65489
rect 116 -65522 208 -65489
rect 614 -65522 706 -65489
rect 581 -65522 614 -65489
rect 738 -65522 830 -65489
rect 240 -65522 332 -65489
rect 830 -65664 863 -65631
rect 332 -65664 365 -65631
rect -9 -65664 83 -65631
rect 83 -65664 116 -65631
rect 116 -65664 208 -65631
rect 738 -65664 830 -65631
rect 240 -65664 332 -65631
rect 489 -65806 581 -65773
rect 830 -65806 863 -65773
rect 365 -65806 457 -65773
rect 332 -65806 365 -65773
rect -9 -65806 83 -65773
rect 83 -65806 116 -65773
rect 116 -65806 208 -65773
rect 614 -65806 706 -65773
rect 581 -65806 614 -65773
rect 738 -65806 830 -65773
rect 489 -65948 581 -65915
rect 830 -65948 863 -65915
rect 365 -65948 457 -65915
rect 332 -65948 365 -65915
rect -9 -65948 83 -65915
rect 83 -65948 116 -65915
rect 116 -65948 208 -65915
rect 614 -65948 706 -65915
rect 581 -65948 614 -65915
rect 738 -65948 830 -65915
rect 863 -65948 955 -65915
rect 830 -66090 863 -66057
rect 365 -66090 457 -66057
rect 332 -66090 365 -66057
rect -9 -66090 83 -66057
rect 83 -66090 116 -66057
rect 116 -66090 208 -66057
rect 614 -66090 706 -66057
rect 581 -66090 614 -66057
rect 738 -66090 830 -66057
rect 863 -66090 955 -66057
rect 830 -66232 863 -66199
rect 489 -66232 581 -66199
rect 332 -66232 365 -66199
rect -9 -66232 83 -66199
rect 83 -66232 116 -66199
rect 116 -66232 208 -66199
rect 614 -66232 706 -66199
rect 365 -66232 457 -66199
rect 738 -66232 830 -66199
rect 581 -66232 614 -66199
rect 489 -66374 581 -66341
rect 830 -66374 863 -66341
rect -9 -66374 83 -66341
rect 83 -66374 116 -66341
rect 116 -66374 208 -66341
rect 581 -66374 614 -66341
rect 738 -66374 830 -66341
rect 863 -66374 955 -66341
rect 830 -66516 863 -66483
rect -9 -66516 83 -66483
rect 83 -66516 116 -66483
rect 116 -66516 208 -66483
rect 614 -66516 706 -66483
rect 581 -66516 614 -66483
rect 738 -66516 830 -66483
rect 830 -66658 863 -66625
rect 489 -66658 581 -66625
rect 365 -66658 457 -66625
rect -9 -66658 83 -66625
rect 332 -66658 365 -66625
rect 83 -66658 116 -66625
rect 116 -66658 208 -66625
rect 614 -66658 706 -66625
rect 581 -66658 614 -66625
rect 738 -66658 830 -66625
rect 240 -66658 332 -66625
rect 863 -66658 955 -66625
rect 489 -66800 581 -66767
rect 830 -66800 863 -66767
rect 365 -66800 457 -66767
rect 332 -66800 365 -66767
rect -9 -66800 83 -66767
rect 83 -66800 116 -66767
rect 614 -66800 706 -66767
rect 581 -66800 614 -66767
rect 240 -66800 332 -66767
rect 863 -66800 955 -66767
rect 830 -66942 863 -66909
rect 365 -66942 457 -66909
rect 332 -66942 365 -66909
rect -9 -66942 83 -66909
rect 83 -66942 116 -66909
rect 614 -66942 706 -66909
rect 581 -66942 614 -66909
rect 738 -66942 830 -66909
rect 240 -66942 332 -66909
rect 863 -66942 955 -66909
rect 830 -67084 863 -67051
rect 489 -67084 581 -67051
rect 332 -67084 365 -67051
rect -9 -67084 83 -67051
rect 83 -67084 116 -67051
rect 614 -67084 706 -67051
rect 365 -67084 457 -67051
rect 581 -67084 614 -67051
rect 240 -67084 332 -67051
rect 863 -67084 955 -67051
rect 489 -67226 581 -67193
rect 830 -67226 863 -67193
rect 332 -67226 365 -67193
rect -9 -67226 83 -67193
rect 83 -67226 116 -67193
rect 614 -67226 706 -67193
rect 581 -67226 614 -67193
rect 738 -67226 830 -67193
rect 240 -67226 332 -67193
rect 863 -67226 955 -67193
rect 830 -67368 863 -67335
rect 332 -67368 365 -67335
rect -9 -67368 83 -67335
rect 83 -67368 116 -67335
rect 614 -67368 706 -67335
rect 581 -67368 614 -67335
rect 738 -67368 830 -67335
rect 240 -67368 332 -67335
rect 863 -67368 955 -67335
rect 489 -67510 581 -67477
rect 830 -67510 863 -67477
rect 365 -67510 457 -67477
rect 332 -67510 365 -67477
rect -9 -67510 83 -67477
rect 83 -67510 116 -67477
rect 614 -67510 706 -67477
rect 581 -67510 614 -67477
rect 738 -67510 830 -67477
rect 863 -67510 955 -67477
rect 489 -67652 581 -67619
rect 830 -67652 863 -67619
rect 365 -67652 457 -67619
rect 332 -67652 365 -67619
rect -9 -67652 83 -67619
rect 83 -67652 116 -67619
rect 614 -67652 706 -67619
rect 581 -67652 614 -67619
rect 863 -67652 955 -67619
rect 830 -67794 863 -67761
rect 489 -67794 581 -67761
rect 332 -67794 365 -67761
rect -9 -67794 83 -67761
rect 83 -67794 116 -67761
rect 614 -67794 706 -67761
rect 365 -67794 457 -67761
rect 738 -67794 830 -67761
rect 581 -67794 614 -67761
rect 863 -67794 955 -67761
rect 489 -67936 581 -67903
rect 830 -67936 863 -67903
rect -9 -67936 83 -67903
rect 83 -67936 116 -67903
rect 614 -67936 706 -67903
rect 581 -67936 614 -67903
rect 863 -67936 955 -67903
rect 830 -68078 863 -68045
rect -9 -68078 83 -68045
rect 83 -68078 116 -68045
rect 614 -68078 706 -68045
rect 581 -68078 614 -68045
rect 738 -68078 830 -68045
rect 863 -68078 955 -68045
rect 489 -68220 581 -68187
rect 365 -68220 457 -68187
rect -9 -68220 83 -68187
rect 332 -68220 365 -68187
rect 83 -68220 116 -68187
rect 116 -68220 208 -68187
rect 614 -68220 706 -68187
rect 581 -68220 614 -68187
rect 240 -68220 332 -68187
rect 489 -68362 581 -68329
rect 830 -68362 863 -68329
rect 365 -68362 457 -68329
rect 332 -68362 365 -68329
rect 83 -68362 116 -68329
rect 116 -68362 208 -68329
rect 614 -68362 706 -68329
rect 581 -68362 614 -68329
rect 738 -68362 830 -68329
rect 240 -68362 332 -68329
rect 863 -68362 955 -68329
rect 830 -68504 863 -68471
rect 332 -68504 365 -68471
rect 83 -68504 116 -68471
rect 116 -68504 208 -68471
rect 365 -68504 457 -68471
rect 738 -68504 830 -68471
rect 240 -68504 332 -68471
rect 863 -68504 955 -68471
rect 489 -68646 581 -68613
rect 830 -68646 863 -68613
rect 332 -68646 365 -68613
rect 83 -68646 116 -68613
rect 116 -68646 208 -68613
rect 614 -68646 706 -68613
rect 581 -68646 614 -68613
rect 738 -68646 830 -68613
rect 240 -68646 332 -68613
rect 863 -68646 955 -68613
rect 830 -68788 863 -68755
rect 332 -68788 365 -68755
rect 83 -68788 116 -68755
rect 116 -68788 208 -68755
rect 614 -68788 706 -68755
rect 581 -68788 614 -68755
rect 738 -68788 830 -68755
rect 240 -68788 332 -68755
rect 863 -68788 955 -68755
rect 830 -68930 863 -68897
rect 489 -68930 581 -68897
rect 365 -68930 457 -68897
rect 332 -68930 365 -68897
rect 83 -68930 116 -68897
rect 116 -68930 208 -68897
rect 614 -68930 706 -68897
rect 581 -68930 614 -68897
rect 240 -68930 332 -68897
rect 863 -68930 955 -68897
rect 489 -69072 581 -69039
rect 830 -69072 863 -69039
rect 365 -69072 457 -69039
rect 332 -69072 365 -69039
rect 83 -69072 116 -69039
rect 116 -69072 208 -69039
rect 581 -69072 614 -69039
rect 738 -69072 830 -69039
rect 830 -69214 863 -69181
rect 365 -69214 457 -69181
rect 332 -69214 365 -69181
rect 83 -69214 116 -69181
rect 116 -69214 208 -69181
rect 614 -69214 706 -69181
rect 581 -69214 614 -69181
rect 738 -69214 830 -69181
rect 863 -69214 955 -69181
rect 830 -69356 863 -69323
rect 489 -69356 581 -69323
rect 83 -69356 116 -69323
rect 116 -69356 208 -69323
rect 614 -69356 706 -69323
rect 581 -69356 614 -69323
rect 738 -69356 830 -69323
rect 863 -69356 955 -69323
rect 489 -69498 581 -69465
rect 830 -69498 863 -69465
rect 83 -69498 116 -69465
rect 116 -69498 208 -69465
rect 614 -69498 706 -69465
rect 581 -69498 614 -69465
rect 738 -69498 830 -69465
rect 863 -69498 955 -69465
rect 830 -69640 863 -69607
rect 83 -69640 116 -69607
rect 116 -69640 208 -69607
rect 738 -69640 830 -69607
rect 863 -69640 955 -69607
rect 489 -69782 581 -69749
rect 830 -69782 863 -69749
rect 365 -69782 457 -69749
rect 332 -69782 365 -69749
rect 614 -69782 706 -69749
rect 581 -69782 614 -69749
rect 738 -69782 830 -69749
rect 240 -69782 332 -69749
rect 863 -69782 955 -69749
rect 489 -69924 581 -69891
rect 830 -69924 863 -69891
rect 365 -69924 457 -69891
rect 332 -69924 365 -69891
rect 614 -69924 706 -69891
rect 581 -69924 614 -69891
rect 738 -69924 830 -69891
rect 240 -69924 332 -69891
rect 863 -69924 955 -69891
rect 830 -70066 863 -70033
rect 365 -70066 457 -70033
rect 332 -70066 365 -70033
rect 614 -70066 706 -70033
rect 581 -70066 614 -70033
rect 240 -70066 332 -70033
rect 863 -70066 955 -70033
rect 830 -70208 863 -70175
rect 489 -70208 581 -70175
rect 332 -70208 365 -70175
rect 614 -70208 706 -70175
rect 581 -70208 614 -70175
rect 738 -70208 830 -70175
rect 240 -70208 332 -70175
rect 863 -70208 955 -70175
rect 489 -70350 581 -70317
rect 830 -70350 863 -70317
rect 332 -70350 365 -70317
rect 581 -70350 614 -70317
rect 738 -70350 830 -70317
rect 240 -70350 332 -70317
rect 830 -70492 863 -70459
rect 332 -70492 365 -70459
rect 614 -70492 706 -70459
rect 581 -70492 614 -70459
rect 738 -70492 830 -70459
rect 240 -70492 332 -70459
rect 863 -70492 955 -70459
rect 830 -70634 863 -70601
rect 489 -70634 581 -70601
rect 365 -70634 457 -70601
rect 332 -70634 365 -70601
rect 614 -70634 706 -70601
rect 581 -70634 614 -70601
rect 738 -70634 830 -70601
rect 240 -70634 332 -70601
rect 863 -70634 955 -70601
rect 489 -70776 581 -70743
rect 830 -70776 863 -70743
rect 365 -70776 457 -70743
rect 332 -70776 365 -70743
rect 614 -70776 706 -70743
rect 581 -70776 614 -70743
rect 738 -70776 830 -70743
rect 863 -70776 955 -70743
rect 489 -70918 581 -70885
rect 830 -70918 863 -70885
rect 365 -70918 457 -70885
rect 332 -70918 365 -70885
rect 614 -70918 706 -70885
rect 581 -70918 614 -70885
rect 738 -70918 830 -70885
rect 863 -70918 955 -70885
rect 830 -71060 863 -71027
rect 365 -71060 457 -71027
rect 332 -71060 365 -71027
rect 614 -71060 706 -71027
rect 581 -71060 614 -71027
rect 863 -71060 955 -71027
rect 830 -71202 863 -71169
rect 332 -71202 365 -71169
rect 365 -71202 457 -71169
rect 738 -71202 830 -71169
rect 863 -71202 955 -71169
rect 830 -71344 863 -71311
rect 489 -71344 581 -71311
rect 614 -71344 706 -71311
rect 581 -71344 614 -71311
rect 738 -71344 830 -71311
rect 863 -71344 955 -71311
rect 830 -71486 863 -71453
rect 489 -71486 581 -71453
rect 614 -71486 706 -71453
rect 581 -71486 614 -71453
rect 738 -71486 830 -71453
rect 863 -71486 955 -71453
rect 489 -71628 581 -71595
rect 830 -71628 863 -71595
rect 581 -71628 614 -71595
rect 738 -71628 830 -71595
rect 863 -71628 955 -71595
rect 830 -71770 863 -71737
rect 614 -71770 706 -71737
rect 581 -71770 614 -71737
rect 738 -71770 830 -71737
rect 863 -71770 955 -71737
rect 581 -71912 614 -71879
rect 614 -71912 706 -71879
rect 830 -71912 863 -71879
rect 863 -71912 955 -71879
rect 830 -72054 863 -72021
rect 614 -72054 706 -72021
rect 581 -72054 614 -72021
rect 738 -72054 830 -72021
rect 863 -72054 955 -72021
rect 738 -72196 830 -72163
rect 830 -72196 863 -72163
rect 830 -72338 863 -72305
rect 863 -72338 955 -72305
rect 830 -72480 863 -72447
rect 863 -72480 955 -72447
rect 904 -9077 955 -9044
rect -9 -9077 42 -9044
rect 655 -9077 706 -9044
rect 489 -9077 540 -9044
rect 406 -9077 457 -9044
rect 240 -9077 291 -9044
rect 157 -9077 208 -9044
rect 738 -9077 789 -9044
rect 904 -9219 955 -9186
rect -9 -9219 42 -9186
rect 655 -9219 706 -9186
rect 489 -9219 540 -9186
rect 406 -9219 457 -9186
rect 240 -9219 291 -9186
rect 157 -9219 208 -9186
rect 738 -9219 789 -9186
rect 904 -9361 955 -9328
rect -9 -9361 42 -9328
rect 655 -9361 706 -9328
rect 489 -9361 540 -9328
rect 406 -9361 457 -9328
rect 240 -9361 291 -9328
rect 157 -9361 208 -9328
rect 738 -9361 789 -9328
rect 904 -9503 955 -9470
rect -9 -9503 42 -9470
rect 655 -9503 706 -9470
rect 489 -9503 540 -9470
rect 406 -9503 457 -9470
rect 240 -9503 291 -9470
rect 157 -9503 208 -9470
rect 738 -9503 789 -9470
rect 904 -9645 955 -9612
rect -9 -9645 42 -9612
rect 655 -9645 706 -9612
rect 489 -9645 540 -9612
rect 406 -9645 457 -9612
rect 240 -9645 291 -9612
rect 157 -9645 208 -9612
rect 738 -9645 789 -9612
rect 904 -9787 955 -9754
rect -9 -9787 42 -9754
rect 655 -9787 706 -9754
rect 489 -9787 540 -9754
rect 406 -9787 457 -9754
rect 240 -9787 291 -9754
rect 157 -9787 208 -9754
rect 738 -9787 789 -9754
rect 904 -9929 955 -9896
rect -9 -9929 42 -9896
rect 655 -9929 706 -9896
rect 489 -9929 540 -9896
rect 406 -9929 457 -9896
rect 240 -9929 291 -9896
rect 157 -9929 208 -9896
rect 738 -9929 789 -9896
rect 904 -10071 955 -10038
rect -9 -10071 42 -10038
rect 655 -10071 706 -10038
rect 489 -10071 540 -10038
rect 406 -10071 457 -10038
rect 240 -10071 291 -10038
rect 157 -10071 208 -10038
rect 738 -10071 789 -10038
rect 904 -10213 955 -10180
rect -9 -10213 42 -10180
rect 655 -10213 706 -10180
rect 489 -10213 540 -10180
rect 406 -10213 457 -10180
rect 240 -10213 291 -10180
rect 157 -10213 208 -10180
rect 738 -10213 789 -10180
rect 904 -10355 955 -10322
rect -9 -10355 42 -10322
rect 655 -10355 706 -10322
rect 489 -10355 540 -10322
rect 406 -10355 457 -10322
rect 240 -10355 291 -10322
rect 157 -10355 208 -10322
rect 738 -10355 789 -10322
rect 904 -10497 955 -10464
rect -9 -10497 42 -10464
rect 655 -10497 706 -10464
rect 489 -10497 540 -10464
rect 406 -10497 457 -10464
rect 240 -10497 291 -10464
rect 157 -10497 208 -10464
rect 738 -10497 789 -10464
rect 904 -10639 955 -10606
rect -9 -10639 42 -10606
rect 655 -10639 706 -10606
rect 489 -10639 540 -10606
rect 406 -10639 457 -10606
rect 240 -10639 291 -10606
rect 157 -10639 208 -10606
rect 738 -10639 789 -10606
rect 904 -10781 955 -10748
rect -9 -10781 42 -10748
rect 655 -10781 706 -10748
rect 489 -10781 540 -10748
rect 406 -10781 457 -10748
rect 240 -10781 291 -10748
rect 157 -10781 208 -10748
rect 738 -10781 789 -10748
rect 904 -10923 955 -10890
rect -9 -10923 42 -10890
rect 655 -10923 706 -10890
rect 489 -10923 540 -10890
rect 406 -10923 457 -10890
rect 240 -10923 291 -10890
rect 157 -10923 208 -10890
rect 738 -10923 789 -10890
rect 904 -11065 955 -11032
rect -9 -11065 42 -11032
rect 655 -11065 706 -11032
rect 489 -11065 540 -11032
rect 406 -11065 457 -11032
rect 240 -11065 291 -11032
rect 157 -11065 208 -11032
rect 738 -11065 789 -11032
rect 904 -11207 955 -11174
rect -9 -11207 42 -11174
rect 655 -11207 706 -11174
rect 489 -11207 540 -11174
rect 406 -11207 457 -11174
rect 240 -11207 291 -11174
rect 157 -11207 208 -11174
rect 738 -11207 789 -11174
rect 904 -11349 955 -11316
rect -9 -11349 42 -11316
rect 655 -11349 706 -11316
rect 489 -11349 540 -11316
rect 406 -11349 457 -11316
rect 240 -11349 291 -11316
rect 157 -11349 208 -11316
rect 738 -11349 789 -11316
rect 904 -11491 955 -11458
rect -9 -11491 42 -11458
rect 655 -11491 706 -11458
rect 489 -11491 540 -11458
rect 406 -11491 457 -11458
rect 240 -11491 291 -11458
rect 157 -11491 208 -11458
rect 738 -11491 789 -11458
rect 904 -11633 955 -11600
rect -9 -11633 42 -11600
rect 655 -11633 706 -11600
rect 489 -11633 540 -11600
rect 406 -11633 457 -11600
rect 240 -11633 291 -11600
rect 157 -11633 208 -11600
rect 738 -11633 789 -11600
rect 904 -11775 955 -11742
rect -9 -11775 42 -11742
rect 655 -11775 706 -11742
rect 489 -11775 540 -11742
rect 406 -11775 457 -11742
rect 240 -11775 291 -11742
rect 157 -11775 208 -11742
rect 738 -11775 789 -11742
rect 904 -11917 955 -11884
rect -9 -11917 42 -11884
rect 655 -11917 706 -11884
rect 489 -11917 540 -11884
rect 406 -11917 457 -11884
rect 240 -11917 291 -11884
rect 157 -11917 208 -11884
rect 738 -11917 789 -11884
rect 904 -12059 955 -12026
rect -9 -12059 42 -12026
rect 655 -12059 706 -12026
rect 489 -12059 540 -12026
rect 406 -12059 457 -12026
rect 240 -12059 291 -12026
rect 157 -12059 208 -12026
rect 738 -12059 789 -12026
rect 904 -12201 955 -12168
rect -9 -12201 42 -12168
rect 655 -12201 706 -12168
rect 489 -12201 540 -12168
rect 406 -12201 457 -12168
rect 240 -12201 291 -12168
rect 157 -12201 208 -12168
rect 738 -12201 789 -12168
rect 904 -12343 955 -12310
rect -9 -12343 42 -12310
rect 655 -12343 706 -12310
rect 489 -12343 540 -12310
rect 406 -12343 457 -12310
rect 240 -12343 291 -12310
rect 157 -12343 208 -12310
rect 738 -12343 789 -12310
rect 904 -12485 955 -12452
rect -9 -12485 42 -12452
rect 655 -12485 706 -12452
rect 489 -12485 540 -12452
rect 406 -12485 457 -12452
rect 240 -12485 291 -12452
rect 157 -12485 208 -12452
rect 738 -12485 789 -12452
rect 904 -12627 955 -12594
rect -9 -12627 42 -12594
rect 655 -12627 706 -12594
rect 489 -12627 540 -12594
rect 406 -12627 457 -12594
rect 240 -12627 291 -12594
rect 157 -12627 208 -12594
rect 738 -12627 789 -12594
rect 904 -12769 955 -12736
rect -9 -12769 42 -12736
rect 655 -12769 706 -12736
rect 489 -12769 540 -12736
rect 406 -12769 457 -12736
rect 240 -12769 291 -12736
rect 157 -12769 208 -12736
rect 738 -12769 789 -12736
rect 904 -12911 955 -12878
rect -9 -12911 42 -12878
rect 655 -12911 706 -12878
rect 489 -12911 540 -12878
rect 406 -12911 457 -12878
rect 240 -12911 291 -12878
rect 157 -12911 208 -12878
rect 738 -12911 789 -12878
rect 904 -13053 955 -13020
rect -9 -13053 42 -13020
rect 655 -13053 706 -13020
rect 489 -13053 540 -13020
rect 406 -13053 457 -13020
rect 240 -13053 291 -13020
rect 157 -13053 208 -13020
rect 738 -13053 789 -13020
rect 904 -13195 955 -13162
rect -9 -13195 42 -13162
rect 655 -13195 706 -13162
rect 489 -13195 540 -13162
rect 406 -13195 457 -13162
rect 240 -13195 291 -13162
rect 157 -13195 208 -13162
rect 738 -13195 789 -13162
rect 904 -13337 955 -13304
rect -9 -13337 42 -13304
rect 655 -13337 706 -13304
rect 489 -13337 540 -13304
rect 406 -13337 457 -13304
rect 240 -13337 291 -13304
rect 157 -13337 208 -13304
rect 738 -13337 789 -13304
rect 904 -13479 955 -13446
rect -9 -13479 42 -13446
rect 655 -13479 706 -13446
rect 489 -13479 540 -13446
rect 406 -13479 457 -13446
rect 240 -13479 291 -13446
rect 157 -13479 208 -13446
rect 738 -13479 789 -13446
rect 904 -13621 955 -13588
rect -9 -13621 42 -13588
rect 655 -13621 706 -13588
rect 489 -13621 540 -13588
rect 406 -13621 457 -13588
rect 240 -13621 291 -13588
rect 157 -13621 208 -13588
rect 738 -13621 789 -13588
rect 904 -13763 955 -13730
rect -9 -13763 42 -13730
rect 655 -13763 706 -13730
rect 489 -13763 540 -13730
rect 406 -13763 457 -13730
rect 240 -13763 291 -13730
rect 157 -13763 208 -13730
rect 738 -13763 789 -13730
rect 904 -13905 955 -13872
rect -9 -13905 42 -13872
rect 655 -13905 706 -13872
rect 489 -13905 540 -13872
rect 406 -13905 457 -13872
rect 240 -13905 291 -13872
rect 157 -13905 208 -13872
rect 738 -13905 789 -13872
rect 904 -14047 955 -14014
rect -9 -14047 42 -14014
rect 655 -14047 706 -14014
rect 489 -14047 540 -14014
rect 406 -14047 457 -14014
rect 240 -14047 291 -14014
rect 157 -14047 208 -14014
rect 738 -14047 789 -14014
rect 904 -14189 955 -14156
rect -9 -14189 42 -14156
rect 655 -14189 706 -14156
rect 489 -14189 540 -14156
rect 406 -14189 457 -14156
rect 240 -14189 291 -14156
rect 157 -14189 208 -14156
rect 738 -14189 789 -14156
rect 904 -14331 955 -14298
rect -9 -14331 42 -14298
rect 655 -14331 706 -14298
rect 489 -14331 540 -14298
rect 406 -14331 457 -14298
rect 240 -14331 291 -14298
rect 157 -14331 208 -14298
rect 738 -14331 789 -14298
rect 904 -14473 955 -14440
rect -9 -14473 42 -14440
rect 655 -14473 706 -14440
rect 489 -14473 540 -14440
rect 406 -14473 457 -14440
rect 240 -14473 291 -14440
rect 157 -14473 208 -14440
rect 738 -14473 789 -14440
rect 904 -14615 955 -14582
rect -9 -14615 42 -14582
rect 655 -14615 706 -14582
rect 489 -14615 540 -14582
rect 406 -14615 457 -14582
rect 240 -14615 291 -14582
rect 157 -14615 208 -14582
rect 738 -14615 789 -14582
rect 904 -14757 955 -14724
rect -9 -14757 42 -14724
rect 655 -14757 706 -14724
rect 489 -14757 540 -14724
rect 406 -14757 457 -14724
rect 240 -14757 291 -14724
rect 157 -14757 208 -14724
rect 738 -14757 789 -14724
rect 904 -14899 955 -14866
rect -9 -14899 42 -14866
rect 655 -14899 706 -14866
rect 489 -14899 540 -14866
rect 406 -14899 457 -14866
rect 240 -14899 291 -14866
rect 157 -14899 208 -14866
rect 738 -14899 789 -14866
rect 904 -15041 955 -15008
rect -9 -15041 42 -15008
rect 655 -15041 706 -15008
rect 489 -15041 540 -15008
rect 406 -15041 457 -15008
rect 240 -15041 291 -15008
rect 157 -15041 208 -15008
rect 738 -15041 789 -15008
rect 904 -15183 955 -15150
rect -9 -15183 42 -15150
rect 655 -15183 706 -15150
rect 489 -15183 540 -15150
rect 406 -15183 457 -15150
rect 240 -15183 291 -15150
rect 157 -15183 208 -15150
rect 738 -15183 789 -15150
rect 904 -15325 955 -15292
rect -9 -15325 42 -15292
rect 655 -15325 706 -15292
rect 489 -15325 540 -15292
rect 406 -15325 457 -15292
rect 240 -15325 291 -15292
rect 157 -15325 208 -15292
rect 738 -15325 789 -15292
rect 904 -15467 955 -15434
rect -9 -15467 42 -15434
rect 655 -15467 706 -15434
rect 489 -15467 540 -15434
rect 406 -15467 457 -15434
rect 240 -15467 291 -15434
rect 157 -15467 208 -15434
rect 738 -15467 789 -15434
rect 904 -15609 955 -15576
rect -9 -15609 42 -15576
rect 655 -15609 706 -15576
rect 489 -15609 540 -15576
rect 406 -15609 457 -15576
rect 240 -15609 291 -15576
rect 157 -15609 208 -15576
rect 738 -15609 789 -15576
rect 904 -15751 955 -15718
rect -9 -15751 42 -15718
rect 655 -15751 706 -15718
rect 489 -15751 540 -15718
rect 406 -15751 457 -15718
rect 240 -15751 291 -15718
rect 157 -15751 208 -15718
rect 738 -15751 789 -15718
rect 904 -15893 955 -15860
rect -9 -15893 42 -15860
rect 655 -15893 706 -15860
rect 489 -15893 540 -15860
rect 406 -15893 457 -15860
rect 240 -15893 291 -15860
rect 157 -15893 208 -15860
rect 738 -15893 789 -15860
rect 904 -16035 955 -16002
rect -9 -16035 42 -16002
rect 655 -16035 706 -16002
rect 489 -16035 540 -16002
rect 406 -16035 457 -16002
rect 240 -16035 291 -16002
rect 157 -16035 208 -16002
rect 738 -16035 789 -16002
rect 904 -16177 955 -16144
rect -9 -16177 42 -16144
rect 655 -16177 706 -16144
rect 489 -16177 540 -16144
rect 406 -16177 457 -16144
rect 240 -16177 291 -16144
rect 157 -16177 208 -16144
rect 738 -16177 789 -16144
rect 904 -16319 955 -16286
rect -9 -16319 42 -16286
rect 655 -16319 706 -16286
rect 489 -16319 540 -16286
rect 406 -16319 457 -16286
rect 240 -16319 291 -16286
rect 157 -16319 208 -16286
rect 738 -16319 789 -16286
rect 904 -16461 955 -16428
rect -9 -16461 42 -16428
rect 655 -16461 706 -16428
rect 489 -16461 540 -16428
rect 406 -16461 457 -16428
rect 240 -16461 291 -16428
rect 157 -16461 208 -16428
rect 738 -16461 789 -16428
rect 904 -16603 955 -16570
rect -9 -16603 42 -16570
rect 655 -16603 706 -16570
rect 489 -16603 540 -16570
rect 406 -16603 457 -16570
rect 240 -16603 291 -16570
rect 157 -16603 208 -16570
rect 738 -16603 789 -16570
rect 904 -16745 955 -16712
rect -9 -16745 42 -16712
rect 655 -16745 706 -16712
rect 489 -16745 540 -16712
rect 406 -16745 457 -16712
rect 240 -16745 291 -16712
rect 157 -16745 208 -16712
rect 738 -16745 789 -16712
rect 904 -16887 955 -16854
rect -9 -16887 42 -16854
rect 655 -16887 706 -16854
rect 489 -16887 540 -16854
rect 406 -16887 457 -16854
rect 240 -16887 291 -16854
rect 157 -16887 208 -16854
rect 738 -16887 789 -16854
rect 904 -17029 955 -16996
rect -9 -17029 42 -16996
rect 655 -17029 706 -16996
rect 489 -17029 540 -16996
rect 406 -17029 457 -16996
rect 240 -17029 291 -16996
rect 157 -17029 208 -16996
rect 738 -17029 789 -16996
rect 904 -17171 955 -17138
rect -9 -17171 42 -17138
rect 655 -17171 706 -17138
rect 489 -17171 540 -17138
rect 406 -17171 457 -17138
rect 240 -17171 291 -17138
rect 157 -17171 208 -17138
rect 738 -17171 789 -17138
rect 904 -17313 955 -17280
rect -9 -17313 42 -17280
rect 655 -17313 706 -17280
rect 489 -17313 540 -17280
rect 406 -17313 457 -17280
rect 240 -17313 291 -17280
rect 157 -17313 208 -17280
rect 738 -17313 789 -17280
rect 904 -17455 955 -17422
rect -9 -17455 42 -17422
rect 655 -17455 706 -17422
rect 489 -17455 540 -17422
rect 406 -17455 457 -17422
rect 240 -17455 291 -17422
rect 157 -17455 208 -17422
rect 738 -17455 789 -17422
rect 904 -17597 955 -17564
rect -9 -17597 42 -17564
rect 655 -17597 706 -17564
rect 489 -17597 540 -17564
rect 406 -17597 457 -17564
rect 240 -17597 291 -17564
rect 157 -17597 208 -17564
rect 738 -17597 789 -17564
rect 904 -17739 955 -17706
rect -9 -17739 42 -17706
rect 655 -17739 706 -17706
rect 489 -17739 540 -17706
rect 406 -17739 457 -17706
rect 240 -17739 291 -17706
rect 157 -17739 208 -17706
rect 738 -17739 789 -17706
rect 904 -17881 955 -17848
rect -9 -17881 42 -17848
rect 655 -17881 706 -17848
rect 489 -17881 540 -17848
rect 406 -17881 457 -17848
rect 240 -17881 291 -17848
rect 157 -17881 208 -17848
rect 738 -17881 789 -17848
rect 904 -18023 955 -17990
rect -9 -18023 42 -17990
rect 655 -18023 706 -17990
rect 489 -18023 540 -17990
rect 406 -18023 457 -17990
rect 240 -18023 291 -17990
rect 157 -18023 208 -17990
rect 738 -18023 789 -17990
rect 904 -18165 955 -18132
rect -9 -18165 42 -18132
rect 655 -18165 706 -18132
rect 489 -18165 540 -18132
rect 406 -18165 457 -18132
rect 240 -18165 291 -18132
rect 157 -18165 208 -18132
rect 738 -18165 789 -18132
rect 738 -18307 789 -18274
rect 904 -18307 955 -18274
rect 904 -18449 955 -18416
rect 655 -18449 706 -18416
rect 738 -18449 789 -18416
rect 904 -18591 955 -18558
rect 489 -18591 540 -18558
rect 738 -18591 789 -18558
rect 904 -18733 955 -18700
rect 655 -18733 706 -18700
rect 489 -18733 540 -18700
rect 738 -18733 789 -18700
rect 904 -18875 955 -18842
rect 406 -18875 457 -18842
rect 738 -18875 789 -18842
rect 904 -19017 955 -18984
rect 406 -19017 457 -18984
rect 655 -19017 706 -18984
rect 738 -19017 789 -18984
rect 904 -19159 955 -19126
rect 406 -19159 457 -19126
rect 489 -19159 540 -19126
rect 738 -19159 789 -19126
rect 904 -19301 955 -19268
rect 655 -19301 706 -19268
rect 489 -19301 540 -19268
rect 406 -19301 457 -19268
rect 738 -19301 789 -19268
rect 904 -19443 955 -19410
rect 240 -19443 291 -19410
rect 738 -19443 789 -19410
rect 904 -19585 955 -19552
rect 655 -19585 706 -19552
rect 240 -19585 291 -19552
rect 738 -19585 789 -19552
rect 904 -19727 955 -19694
rect 489 -19727 540 -19694
rect 240 -19727 291 -19694
rect 738 -19727 789 -19694
rect 904 -19869 955 -19836
rect 655 -19869 706 -19836
rect 489 -19869 540 -19836
rect 240 -19869 291 -19836
rect 738 -19869 789 -19836
rect 904 -20011 955 -19978
rect 406 -20011 457 -19978
rect 240 -20011 291 -19978
rect 738 -20011 789 -19978
rect 904 -20153 955 -20120
rect 406 -20153 457 -20120
rect 655 -20153 706 -20120
rect 240 -20153 291 -20120
rect 738 -20153 789 -20120
rect 904 -20295 955 -20262
rect 406 -20295 457 -20262
rect 489 -20295 540 -20262
rect 240 -20295 291 -20262
rect 738 -20295 789 -20262
rect 904 -20437 955 -20404
rect 655 -20437 706 -20404
rect 489 -20437 540 -20404
rect 406 -20437 457 -20404
rect 240 -20437 291 -20404
rect 738 -20437 789 -20404
rect 904 -20579 955 -20546
rect 157 -20579 208 -20546
rect 738 -20579 789 -20546
rect 904 -20721 955 -20688
rect 655 -20721 706 -20688
rect 157 -20721 208 -20688
rect 738 -20721 789 -20688
rect 904 -20863 955 -20830
rect 489 -20863 540 -20830
rect 157 -20863 208 -20830
rect 738 -20863 789 -20830
rect 904 -21005 955 -20972
rect 655 -21005 706 -20972
rect 489 -21005 540 -20972
rect 157 -21005 208 -20972
rect 738 -21005 789 -20972
rect 904 -21147 955 -21114
rect 406 -21147 457 -21114
rect 157 -21147 208 -21114
rect 738 -21147 789 -21114
rect 904 -21289 955 -21256
rect 406 -21289 457 -21256
rect 655 -21289 706 -21256
rect 157 -21289 208 -21256
rect 738 -21289 789 -21256
rect 904 -21431 955 -21398
rect 406 -21431 457 -21398
rect 489 -21431 540 -21398
rect 157 -21431 208 -21398
rect 738 -21431 789 -21398
rect 904 -21573 955 -21540
rect 655 -21573 706 -21540
rect 489 -21573 540 -21540
rect 406 -21573 457 -21540
rect 157 -21573 208 -21540
rect 738 -21573 789 -21540
rect 904 -21715 955 -21682
rect 240 -21715 291 -21682
rect 157 -21715 208 -21682
rect 738 -21715 789 -21682
rect 904 -21857 955 -21824
rect 655 -21857 706 -21824
rect 240 -21857 291 -21824
rect 157 -21857 208 -21824
rect 738 -21857 789 -21824
rect 904 -21999 955 -21966
rect 489 -21999 540 -21966
rect 240 -21999 291 -21966
rect 157 -21999 208 -21966
rect 738 -21999 789 -21966
rect 904 -22141 955 -22108
rect 655 -22141 706 -22108
rect 489 -22141 540 -22108
rect 240 -22141 291 -22108
rect 157 -22141 208 -22108
rect 738 -22141 789 -22108
rect 904 -22283 955 -22250
rect 406 -22283 457 -22250
rect 240 -22283 291 -22250
rect 157 -22283 208 -22250
rect 738 -22283 789 -22250
rect 904 -22425 955 -22392
rect 406 -22425 457 -22392
rect 655 -22425 706 -22392
rect 240 -22425 291 -22392
rect 157 -22425 208 -22392
rect 738 -22425 789 -22392
rect 904 -22567 955 -22534
rect 406 -22567 457 -22534
rect 489 -22567 540 -22534
rect 240 -22567 291 -22534
rect 157 -22567 208 -22534
rect 738 -22567 789 -22534
rect 904 -22709 955 -22676
rect 655 -22709 706 -22676
rect 489 -22709 540 -22676
rect 406 -22709 457 -22676
rect 240 -22709 291 -22676
rect 157 -22709 208 -22676
rect 738 -22709 789 -22676
rect 904 -22851 955 -22818
rect -9 -22851 42 -22818
rect 738 -22851 789 -22818
rect 904 -22993 955 -22960
rect -9 -22993 42 -22960
rect 655 -22993 706 -22960
rect 738 -22993 789 -22960
rect 904 -23135 955 -23102
rect -9 -23135 42 -23102
rect 489 -23135 540 -23102
rect 738 -23135 789 -23102
rect 904 -23277 955 -23244
rect -9 -23277 42 -23244
rect 655 -23277 706 -23244
rect 489 -23277 540 -23244
rect 738 -23277 789 -23244
rect 904 -23419 955 -23386
rect -9 -23419 42 -23386
rect 406 -23419 457 -23386
rect 738 -23419 789 -23386
rect 904 -23561 955 -23528
rect -9 -23561 42 -23528
rect 406 -23561 457 -23528
rect 655 -23561 706 -23528
rect 738 -23561 789 -23528
rect 904 -23703 955 -23670
rect -9 -23703 42 -23670
rect 406 -23703 457 -23670
rect 489 -23703 540 -23670
rect 738 -23703 789 -23670
rect 904 -23845 955 -23812
rect -9 -23845 42 -23812
rect 655 -23845 706 -23812
rect 489 -23845 540 -23812
rect 406 -23845 457 -23812
rect 738 -23845 789 -23812
rect 904 -23987 955 -23954
rect -9 -23987 42 -23954
rect 240 -23987 291 -23954
rect 738 -23987 789 -23954
rect 904 -24129 955 -24096
rect -9 -24129 42 -24096
rect 655 -24129 706 -24096
rect 240 -24129 291 -24096
rect 738 -24129 789 -24096
rect 904 -24271 955 -24238
rect -9 -24271 42 -24238
rect 489 -24271 540 -24238
rect 240 -24271 291 -24238
rect 738 -24271 789 -24238
rect 904 -24413 955 -24380
rect -9 -24413 42 -24380
rect 655 -24413 706 -24380
rect 489 -24413 540 -24380
rect 240 -24413 291 -24380
rect 738 -24413 789 -24380
rect 904 -24555 955 -24522
rect -9 -24555 42 -24522
rect 406 -24555 457 -24522
rect 240 -24555 291 -24522
rect 738 -24555 789 -24522
rect 904 -24697 955 -24664
rect -9 -24697 42 -24664
rect 406 -24697 457 -24664
rect 655 -24697 706 -24664
rect 240 -24697 291 -24664
rect 738 -24697 789 -24664
rect 904 -24839 955 -24806
rect -9 -24839 42 -24806
rect 406 -24839 457 -24806
rect 489 -24839 540 -24806
rect 240 -24839 291 -24806
rect 738 -24839 789 -24806
rect 904 -24981 955 -24948
rect -9 -24981 42 -24948
rect 655 -24981 706 -24948
rect 489 -24981 540 -24948
rect 406 -24981 457 -24948
rect 240 -24981 291 -24948
rect 738 -24981 789 -24948
rect 904 -25123 955 -25090
rect -9 -25123 42 -25090
rect 157 -25123 208 -25090
rect 738 -25123 789 -25090
rect 904 -25265 955 -25232
rect -9 -25265 42 -25232
rect 655 -25265 706 -25232
rect 157 -25265 208 -25232
rect 738 -25265 789 -25232
rect 904 -25407 955 -25374
rect -9 -25407 42 -25374
rect 489 -25407 540 -25374
rect 157 -25407 208 -25374
rect 738 -25407 789 -25374
rect 904 -25549 955 -25516
rect -9 -25549 42 -25516
rect 655 -25549 706 -25516
rect 489 -25549 540 -25516
rect 157 -25549 208 -25516
rect 738 -25549 789 -25516
rect 904 -25691 955 -25658
rect -9 -25691 42 -25658
rect 406 -25691 457 -25658
rect 157 -25691 208 -25658
rect 738 -25691 789 -25658
rect 904 -25833 955 -25800
rect -9 -25833 42 -25800
rect 406 -25833 457 -25800
rect 655 -25833 706 -25800
rect 157 -25833 208 -25800
rect 738 -25833 789 -25800
rect 904 -25975 955 -25942
rect -9 -25975 42 -25942
rect 406 -25975 457 -25942
rect 489 -25975 540 -25942
rect 157 -25975 208 -25942
rect 738 -25975 789 -25942
rect 904 -26117 955 -26084
rect -9 -26117 42 -26084
rect 655 -26117 706 -26084
rect 489 -26117 540 -26084
rect 406 -26117 457 -26084
rect 157 -26117 208 -26084
rect 738 -26117 789 -26084
rect 904 -26259 955 -26226
rect -9 -26259 42 -26226
rect 240 -26259 291 -26226
rect 157 -26259 208 -26226
rect 738 -26259 789 -26226
rect 904 -26401 955 -26368
rect -9 -26401 42 -26368
rect 655 -26401 706 -26368
rect 240 -26401 291 -26368
rect 157 -26401 208 -26368
rect 738 -26401 789 -26368
rect 904 -26543 955 -26510
rect -9 -26543 42 -26510
rect 489 -26543 540 -26510
rect 240 -26543 291 -26510
rect 157 -26543 208 -26510
rect 738 -26543 789 -26510
rect 904 -26685 955 -26652
rect -9 -26685 42 -26652
rect 655 -26685 706 -26652
rect 489 -26685 540 -26652
rect 240 -26685 291 -26652
rect 157 -26685 208 -26652
rect 738 -26685 789 -26652
rect 904 -26827 955 -26794
rect -9 -26827 42 -26794
rect 406 -26827 457 -26794
rect 240 -26827 291 -26794
rect 157 -26827 208 -26794
rect 738 -26827 789 -26794
rect 904 -26969 955 -26936
rect -9 -26969 42 -26936
rect 406 -26969 457 -26936
rect 655 -26969 706 -26936
rect 240 -26969 291 -26936
rect 157 -26969 208 -26936
rect 738 -26969 789 -26936
rect 904 -27111 955 -27078
rect -9 -27111 42 -27078
rect 406 -27111 457 -27078
rect 489 -27111 540 -27078
rect 240 -27111 291 -27078
rect 157 -27111 208 -27078
rect 738 -27111 789 -27078
rect 904 -27253 955 -27220
rect -9 -27253 42 -27220
rect 655 -27253 706 -27220
rect 489 -27253 540 -27220
rect 406 -27253 457 -27220
rect 240 -27253 291 -27220
rect 157 -27253 208 -27220
rect 738 -27253 789 -27220
rect 904 -27395 955 -27362
rect -9 -27395 42 -27362
rect 655 -27395 706 -27362
rect 489 -27395 540 -27362
rect 406 -27395 457 -27362
rect 240 -27395 291 -27362
rect 157 -27395 208 -27362
rect 738 -27395 789 -27362
rect 904 -27537 955 -27504
rect -9 -27537 42 -27504
rect 406 -27537 457 -27504
rect 489 -27537 540 -27504
rect 240 -27537 291 -27504
rect 157 -27537 208 -27504
rect 738 -27537 789 -27504
rect 655 -27537 706 -27504
rect 904 -27679 955 -27646
rect -9 -27679 42 -27646
rect 406 -27679 457 -27646
rect 655 -27679 706 -27646
rect 240 -27679 291 -27646
rect 157 -27679 208 -27646
rect 738 -27679 789 -27646
rect 904 -27821 955 -27788
rect -9 -27821 42 -27788
rect 406 -27821 457 -27788
rect 655 -27821 706 -27788
rect 240 -27821 291 -27788
rect 157 -27821 208 -27788
rect 738 -27821 789 -27788
rect 489 -27821 540 -27788
rect 904 -27963 955 -27930
rect -9 -27963 42 -27930
rect 655 -27963 706 -27930
rect 489 -27963 540 -27930
rect 240 -27963 291 -27930
rect 157 -27963 208 -27930
rect 738 -27963 789 -27930
rect 904 -28105 955 -28072
rect -9 -28105 42 -28072
rect 489 -28105 540 -28072
rect 655 -28105 706 -28072
rect 240 -28105 291 -28072
rect 157 -28105 208 -28072
rect 738 -28105 789 -28072
rect 904 -28247 955 -28214
rect -9 -28247 42 -28214
rect 655 -28247 706 -28214
rect 240 -28247 291 -28214
rect 157 -28247 208 -28214
rect 738 -28247 789 -28214
rect 904 -28389 955 -28356
rect -9 -28389 42 -28356
rect 655 -28389 706 -28356
rect 489 -28389 540 -28356
rect 240 -28389 291 -28356
rect 157 -28389 208 -28356
rect 738 -28389 789 -28356
rect 406 -28389 457 -28356
rect 904 -28531 955 -28498
rect -9 -28531 42 -28498
rect 655 -28531 706 -28498
rect 489 -28531 540 -28498
rect 406 -28531 457 -28498
rect 157 -28531 208 -28498
rect 738 -28531 789 -28498
rect 904 -28673 955 -28640
rect -9 -28673 42 -28640
rect 406 -28673 457 -28640
rect 489 -28673 540 -28640
rect 655 -28673 706 -28640
rect 157 -28673 208 -28640
rect 738 -28673 789 -28640
rect 904 -28815 955 -28782
rect -9 -28815 42 -28782
rect 406 -28815 457 -28782
rect 655 -28815 706 -28782
rect 157 -28815 208 -28782
rect 738 -28815 789 -28782
rect 904 -28957 955 -28924
rect -9 -28957 42 -28924
rect 406 -28957 457 -28924
rect 655 -28957 706 -28924
rect 489 -28957 540 -28924
rect 157 -28957 208 -28924
rect 738 -28957 789 -28924
rect 904 -29099 955 -29066
rect -9 -29099 42 -29066
rect 655 -29099 706 -29066
rect 489 -29099 540 -29066
rect 157 -29099 208 -29066
rect 738 -29099 789 -29066
rect 904 -29241 955 -29208
rect -9 -29241 42 -29208
rect 489 -29241 540 -29208
rect 655 -29241 706 -29208
rect 157 -29241 208 -29208
rect 738 -29241 789 -29208
rect 904 -29383 955 -29350
rect -9 -29383 42 -29350
rect 655 -29383 706 -29350
rect 157 -29383 208 -29350
rect 738 -29383 789 -29350
rect 904 -29525 955 -29492
rect 240 -29525 291 -29492
rect -9 -29525 42 -29492
rect 655 -29525 706 -29492
rect 489 -29525 540 -29492
rect 406 -29525 457 -29492
rect 157 -29525 208 -29492
rect 738 -29525 789 -29492
rect 904 -29667 955 -29634
rect -9 -29667 42 -29634
rect 655 -29667 706 -29634
rect 489 -29667 540 -29634
rect 406 -29667 457 -29634
rect 240 -29667 291 -29634
rect 738 -29667 789 -29634
rect 904 -29809 955 -29776
rect -9 -29809 42 -29776
rect 406 -29809 457 -29776
rect 489 -29809 540 -29776
rect 655 -29809 706 -29776
rect 240 -29809 291 -29776
rect 738 -29809 789 -29776
rect 904 -29951 955 -29918
rect -9 -29951 42 -29918
rect 406 -29951 457 -29918
rect 655 -29951 706 -29918
rect 240 -29951 291 -29918
rect 738 -29951 789 -29918
rect 904 -30093 955 -30060
rect -9 -30093 42 -30060
rect 406 -30093 457 -30060
rect 655 -30093 706 -30060
rect 240 -30093 291 -30060
rect 489 -30093 540 -30060
rect 738 -30093 789 -30060
rect 904 -30235 955 -30202
rect -9 -30235 42 -30202
rect 655 -30235 706 -30202
rect 489 -30235 540 -30202
rect 240 -30235 291 -30202
rect 738 -30235 789 -30202
rect 904 -30377 955 -30344
rect -9 -30377 42 -30344
rect 655 -30377 706 -30344
rect 489 -30377 540 -30344
rect 240 -30377 291 -30344
rect 738 -30377 789 -30344
rect 904 -30519 955 -30486
rect -9 -30519 42 -30486
rect 655 -30519 706 -30486
rect 240 -30519 291 -30486
rect 738 -30519 789 -30486
rect 904 -30661 955 -30628
rect -9 -30661 42 -30628
rect 655 -30661 706 -30628
rect 489 -30661 540 -30628
rect 406 -30661 457 -30628
rect 240 -30661 291 -30628
rect 738 -30661 789 -30628
rect 904 -30803 955 -30770
rect -9 -30803 42 -30770
rect 655 -30803 706 -30770
rect 489 -30803 540 -30770
rect 406 -30803 457 -30770
rect 738 -30803 789 -30770
rect 904 -30945 955 -30912
rect -9 -30945 42 -30912
rect 406 -30945 457 -30912
rect 489 -30945 540 -30912
rect 655 -30945 706 -30912
rect 738 -30945 789 -30912
rect 904 -31087 955 -31054
rect -9 -31087 42 -31054
rect 406 -31087 457 -31054
rect 655 -31087 706 -31054
rect 738 -31087 789 -31054
rect 904 -31229 955 -31196
rect -9 -31229 42 -31196
rect 406 -31229 457 -31196
rect 655 -31229 706 -31196
rect 489 -31229 540 -31196
rect 738 -31229 789 -31196
rect 904 -31371 955 -31338
rect -9 -31371 42 -31338
rect 655 -31371 706 -31338
rect 489 -31371 540 -31338
rect 738 -31371 789 -31338
rect 904 -31513 955 -31480
rect -9 -31513 42 -31480
rect 655 -31513 706 -31480
rect 489 -31513 540 -31480
rect 738 -31513 789 -31480
rect 904 -31655 955 -31622
rect -9 -31655 42 -31622
rect 655 -31655 706 -31622
rect 738 -31655 789 -31622
rect 904 -31797 955 -31764
rect -9 -31797 42 -31764
rect 655 -31797 706 -31764
rect 489 -31797 540 -31764
rect 406 -31797 457 -31764
rect 240 -31797 291 -31764
rect 157 -31797 208 -31764
rect 738 -31797 789 -31764
rect 904 -31939 955 -31906
rect 655 -31939 706 -31906
rect 489 -31939 540 -31906
rect 406 -31939 457 -31906
rect 240 -31939 291 -31906
rect 157 -31939 208 -31906
rect 738 -31939 789 -31906
rect 904 -32081 955 -32048
rect 406 -32081 457 -32048
rect 489 -32081 540 -32048
rect 240 -32081 291 -32048
rect 157 -32081 208 -32048
rect 738 -32081 789 -32048
rect 655 -32081 706 -32048
rect 904 -32223 955 -32190
rect 406 -32223 457 -32190
rect 655 -32223 706 -32190
rect 240 -32223 291 -32190
rect 157 -32223 208 -32190
rect 738 -32223 789 -32190
rect 904 -32365 955 -32332
rect 406 -32365 457 -32332
rect 655 -32365 706 -32332
rect 240 -32365 291 -32332
rect 157 -32365 208 -32332
rect 738 -32365 789 -32332
rect 489 -32365 540 -32332
rect 904 -32507 955 -32474
rect 655 -32507 706 -32474
rect 489 -32507 540 -32474
rect 240 -32507 291 -32474
rect 157 -32507 208 -32474
rect 738 -32507 789 -32474
rect 904 -32649 955 -32616
rect 489 -32649 540 -32616
rect 655 -32649 706 -32616
rect 240 -32649 291 -32616
rect 157 -32649 208 -32616
rect 738 -32649 789 -32616
rect 904 -32791 955 -32758
rect 655 -32791 706 -32758
rect 240 -32791 291 -32758
rect 157 -32791 208 -32758
rect 738 -32791 789 -32758
rect 904 -32933 955 -32900
rect 655 -32933 706 -32900
rect 489 -32933 540 -32900
rect 240 -32933 291 -32900
rect 157 -32933 208 -32900
rect 738 -32933 789 -32900
rect 406 -32933 457 -32900
rect 904 -33075 955 -33042
rect 655 -33075 706 -33042
rect 489 -33075 540 -33042
rect 406 -33075 457 -33042
rect 157 -33075 208 -33042
rect 738 -33075 789 -33042
rect 904 -33217 955 -33184
rect 406 -33217 457 -33184
rect 489 -33217 540 -33184
rect 655 -33217 706 -33184
rect 157 -33217 208 -33184
rect 738 -33217 789 -33184
rect 904 -33359 955 -33326
rect 406 -33359 457 -33326
rect 655 -33359 706 -33326
rect 157 -33359 208 -33326
rect 738 -33359 789 -33326
rect 904 -33501 955 -33468
rect 406 -33501 457 -33468
rect 655 -33501 706 -33468
rect 489 -33501 540 -33468
rect 157 -33501 208 -33468
rect 738 -33501 789 -33468
rect 904 -33643 955 -33610
rect 655 -33643 706 -33610
rect 489 -33643 540 -33610
rect 157 -33643 208 -33610
rect 738 -33643 789 -33610
rect 904 -33785 955 -33752
rect 489 -33785 540 -33752
rect 655 -33785 706 -33752
rect 157 -33785 208 -33752
rect 738 -33785 789 -33752
rect 904 -33927 955 -33894
rect 655 -33927 706 -33894
rect 157 -33927 208 -33894
rect 738 -33927 789 -33894
rect 904 -34069 955 -34036
rect 240 -34069 291 -34036
rect 655 -34069 706 -34036
rect 489 -34069 540 -34036
rect 406 -34069 457 -34036
rect 157 -34069 208 -34036
rect 738 -34069 789 -34036
rect 904 -34211 955 -34178
rect 655 -34211 706 -34178
rect 489 -34211 540 -34178
rect 406 -34211 457 -34178
rect 240 -34211 291 -34178
rect 738 -34211 789 -34178
rect 904 -34353 955 -34320
rect 406 -34353 457 -34320
rect 489 -34353 540 -34320
rect 655 -34353 706 -34320
rect 240 -34353 291 -34320
rect 738 -34353 789 -34320
rect 904 -34495 955 -34462
rect 406 -34495 457 -34462
rect 655 -34495 706 -34462
rect 240 -34495 291 -34462
rect 738 -34495 789 -34462
rect 904 -34637 955 -34604
rect 406 -34637 457 -34604
rect 655 -34637 706 -34604
rect 240 -34637 291 -34604
rect 489 -34637 540 -34604
rect 738 -34637 789 -34604
rect 904 -34779 955 -34746
rect 655 -34779 706 -34746
rect 489 -34779 540 -34746
rect 240 -34779 291 -34746
rect 738 -34779 789 -34746
rect 904 -34921 955 -34888
rect 655 -34921 706 -34888
rect 489 -34921 540 -34888
rect 240 -34921 291 -34888
rect 738 -34921 789 -34888
rect 904 -35063 955 -35030
rect 655 -35063 706 -35030
rect 240 -35063 291 -35030
rect 738 -35063 789 -35030
rect 904 -35205 955 -35172
rect 655 -35205 706 -35172
rect 489 -35205 540 -35172
rect 406 -35205 457 -35172
rect 240 -35205 291 -35172
rect 738 -35205 789 -35172
rect 904 -35347 955 -35314
rect 655 -35347 706 -35314
rect 489 -35347 540 -35314
rect 406 -35347 457 -35314
rect 738 -35347 789 -35314
rect 904 -35489 955 -35456
rect 406 -35489 457 -35456
rect 489 -35489 540 -35456
rect 655 -35489 706 -35456
rect 738 -35489 789 -35456
rect 904 -35631 955 -35598
rect 406 -35631 457 -35598
rect 655 -35631 706 -35598
rect 738 -35631 789 -35598
rect 904 -35773 955 -35740
rect 406 -35773 457 -35740
rect 655 -35773 706 -35740
rect 489 -35773 540 -35740
rect 738 -35773 789 -35740
rect 904 -35915 955 -35882
rect 655 -35915 706 -35882
rect 489 -35915 540 -35882
rect 738 -35915 789 -35882
rect 904 -36057 955 -36024
rect 655 -36057 706 -36024
rect 489 -36057 540 -36024
rect 738 -36057 789 -36024
rect 904 -36199 955 -36166
rect 655 -36199 706 -36166
rect 738 -36199 789 -36166
rect 904 -36341 955 -36308
rect 904 -36483 955 -36450
rect 904 -36625 955 -36592
rect 738 -36625 789 -36592
rect 904 -36767 955 -36734
rect 655 -36767 706 -36734
rect 904 -36909 955 -36876
rect 655 -36909 706 -36876
rect 738 -36909 789 -36876
rect 904 -37051 955 -37018
rect 489 -37051 540 -37018
rect 904 -37193 955 -37160
rect 489 -37193 540 -37160
rect 738 -37193 789 -37160
rect 904 -37335 955 -37302
rect 655 -37335 706 -37302
rect 489 -37335 540 -37302
rect 904 -37477 955 -37444
rect 655 -37477 706 -37444
rect 489 -37477 540 -37444
rect 738 -37477 789 -37444
rect 904 -37619 955 -37586
rect 406 -37619 457 -37586
rect 904 -37761 955 -37728
rect 406 -37761 457 -37728
rect 738 -37761 789 -37728
rect 904 -37903 955 -37870
rect 406 -37903 457 -37870
rect 655 -37903 706 -37870
rect 904 -38045 955 -38012
rect 655 -38045 706 -38012
rect 406 -38045 457 -38012
rect 738 -38045 789 -38012
rect 904 -38187 955 -38154
rect 406 -38187 457 -38154
rect 489 -38187 540 -38154
rect 904 -38329 955 -38296
rect 406 -38329 457 -38296
rect 489 -38329 540 -38296
rect 738 -38329 789 -38296
rect 904 -38471 955 -38438
rect 406 -38471 457 -38438
rect 655 -38471 706 -38438
rect 489 -38471 540 -38438
rect 904 -38613 955 -38580
rect 655 -38613 706 -38580
rect 489 -38613 540 -38580
rect 406 -38613 457 -38580
rect 738 -38613 789 -38580
rect 240 -38755 291 -38722
rect 904 -38755 955 -38722
rect 904 -38897 955 -38864
rect 240 -38897 291 -38864
rect 738 -38897 789 -38864
rect 904 -39039 955 -39006
rect 655 -39039 706 -39006
rect 240 -39039 291 -39006
rect 904 -39181 955 -39148
rect 655 -39181 706 -39148
rect 240 -39181 291 -39148
rect 738 -39181 789 -39148
rect 904 -39323 955 -39290
rect 489 -39323 540 -39290
rect 240 -39323 291 -39290
rect 904 -39465 955 -39432
rect 489 -39465 540 -39432
rect 240 -39465 291 -39432
rect 738 -39465 789 -39432
rect 904 -39607 955 -39574
rect 655 -39607 706 -39574
rect 489 -39607 540 -39574
rect 240 -39607 291 -39574
rect 904 -39749 955 -39716
rect 655 -39749 706 -39716
rect 489 -39749 540 -39716
rect 240 -39749 291 -39716
rect 738 -39749 789 -39716
rect 904 -39891 955 -39858
rect 406 -39891 457 -39858
rect 240 -39891 291 -39858
rect 904 -40033 955 -40000
rect 406 -40033 457 -40000
rect 240 -40033 291 -40000
rect 738 -40033 789 -40000
rect 904 -40175 955 -40142
rect 406 -40175 457 -40142
rect 655 -40175 706 -40142
rect 240 -40175 291 -40142
rect 904 -40317 955 -40284
rect 655 -40317 706 -40284
rect 406 -40317 457 -40284
rect 240 -40317 291 -40284
rect 738 -40317 789 -40284
rect 904 -40459 955 -40426
rect 406 -40459 457 -40426
rect 489 -40459 540 -40426
rect 240 -40459 291 -40426
rect 904 -40601 955 -40568
rect 406 -40601 457 -40568
rect 489 -40601 540 -40568
rect 240 -40601 291 -40568
rect 738 -40601 789 -40568
rect 904 -40743 955 -40710
rect 406 -40743 457 -40710
rect 655 -40743 706 -40710
rect 489 -40743 540 -40710
rect 240 -40743 291 -40710
rect 904 -40885 955 -40852
rect 655 -40885 706 -40852
rect 489 -40885 540 -40852
rect 406 -40885 457 -40852
rect 240 -40885 291 -40852
rect 738 -40885 789 -40852
rect 157 -41027 208 -40994
rect 904 -41027 955 -40994
rect 904 -41169 955 -41136
rect 157 -41169 208 -41136
rect 738 -41169 789 -41136
rect 904 -41311 955 -41278
rect 655 -41311 706 -41278
rect 157 -41311 208 -41278
rect 904 -41453 955 -41420
rect 655 -41453 706 -41420
rect 157 -41453 208 -41420
rect 738 -41453 789 -41420
rect 904 -41595 955 -41562
rect 489 -41595 540 -41562
rect 157 -41595 208 -41562
rect 904 -41737 955 -41704
rect 489 -41737 540 -41704
rect 157 -41737 208 -41704
rect 738 -41737 789 -41704
rect 904 -41879 955 -41846
rect 655 -41879 706 -41846
rect 489 -41879 540 -41846
rect 157 -41879 208 -41846
rect 904 -42021 955 -41988
rect 655 -42021 706 -41988
rect 489 -42021 540 -41988
rect 157 -42021 208 -41988
rect 738 -42021 789 -41988
rect 904 -42163 955 -42130
rect 406 -42163 457 -42130
rect 157 -42163 208 -42130
rect 904 -42305 955 -42272
rect 406 -42305 457 -42272
rect 157 -42305 208 -42272
rect 738 -42305 789 -42272
rect 904 -42447 955 -42414
rect 406 -42447 457 -42414
rect 655 -42447 706 -42414
rect 157 -42447 208 -42414
rect 904 -42589 955 -42556
rect 655 -42589 706 -42556
rect 406 -42589 457 -42556
rect 157 -42589 208 -42556
rect 738 -42589 789 -42556
rect 904 -42731 955 -42698
rect 406 -42731 457 -42698
rect 489 -42731 540 -42698
rect 157 -42731 208 -42698
rect 904 -42873 955 -42840
rect 406 -42873 457 -42840
rect 489 -42873 540 -42840
rect 157 -42873 208 -42840
rect 738 -42873 789 -42840
rect 904 -43015 955 -42982
rect 406 -43015 457 -42982
rect 655 -43015 706 -42982
rect 489 -43015 540 -42982
rect 157 -43015 208 -42982
rect 904 -43157 955 -43124
rect 655 -43157 706 -43124
rect 489 -43157 540 -43124
rect 406 -43157 457 -43124
rect 157 -43157 208 -43124
rect 738 -43157 789 -43124
rect 904 -43299 955 -43266
rect 240 -43299 291 -43266
rect 157 -43299 208 -43266
rect 904 -43441 955 -43408
rect 240 -43441 291 -43408
rect 157 -43441 208 -43408
rect 738 -43441 789 -43408
rect 904 -43583 955 -43550
rect 655 -43583 706 -43550
rect 240 -43583 291 -43550
rect 157 -43583 208 -43550
rect 904 -43725 955 -43692
rect 655 -43725 706 -43692
rect 240 -43725 291 -43692
rect 157 -43725 208 -43692
rect 738 -43725 789 -43692
rect 904 -43867 955 -43834
rect 489 -43867 540 -43834
rect 240 -43867 291 -43834
rect 157 -43867 208 -43834
rect 904 -44009 955 -43976
rect 489 -44009 540 -43976
rect 240 -44009 291 -43976
rect 157 -44009 208 -43976
rect 738 -44009 789 -43976
rect 904 -44151 955 -44118
rect 655 -44151 706 -44118
rect 489 -44151 540 -44118
rect 240 -44151 291 -44118
rect 157 -44151 208 -44118
rect 904 -44293 955 -44260
rect 655 -44293 706 -44260
rect 489 -44293 540 -44260
rect 240 -44293 291 -44260
rect 157 -44293 208 -44260
rect 738 -44293 789 -44260
rect 904 -44435 955 -44402
rect 406 -44435 457 -44402
rect 240 -44435 291 -44402
rect 157 -44435 208 -44402
rect 904 -44577 955 -44544
rect 406 -44577 457 -44544
rect 240 -44577 291 -44544
rect 157 -44577 208 -44544
rect 738 -44577 789 -44544
rect 904 -44719 955 -44686
rect 406 -44719 457 -44686
rect 655 -44719 706 -44686
rect 240 -44719 291 -44686
rect 157 -44719 208 -44686
rect 904 -44861 955 -44828
rect 655 -44861 706 -44828
rect 406 -44861 457 -44828
rect 240 -44861 291 -44828
rect 157 -44861 208 -44828
rect 738 -44861 789 -44828
rect 904 -45003 955 -44970
rect 406 -45003 457 -44970
rect 489 -45003 540 -44970
rect 240 -45003 291 -44970
rect 157 -45003 208 -44970
rect 904 -45145 955 -45112
rect 406 -45145 457 -45112
rect 489 -45145 540 -45112
rect 240 -45145 291 -45112
rect 157 -45145 208 -45112
rect 738 -45145 789 -45112
rect 904 -45287 955 -45254
rect 406 -45287 457 -45254
rect 655 -45287 706 -45254
rect 489 -45287 540 -45254
rect 240 -45287 291 -45254
rect 157 -45287 208 -45254
rect 904 -45429 955 -45396
rect 655 -45429 706 -45396
rect 489 -45429 540 -45396
rect 406 -45429 457 -45396
rect 240 -45429 291 -45396
rect 157 -45429 208 -45396
rect 738 -45429 789 -45396
rect -9 -45571 42 -45538
rect 904 -45571 955 -45538
rect 904 -45713 955 -45680
rect -9 -45713 42 -45680
rect 738 -45713 789 -45680
rect 904 -45855 955 -45822
rect -9 -45855 42 -45822
rect 655 -45855 706 -45822
rect 904 -45997 955 -45964
rect -9 -45997 42 -45964
rect 655 -45997 706 -45964
rect 738 -45997 789 -45964
rect 904 -46139 955 -46106
rect -9 -46139 42 -46106
rect 489 -46139 540 -46106
rect 904 -46281 955 -46248
rect -9 -46281 42 -46248
rect 489 -46281 540 -46248
rect 738 -46281 789 -46248
rect 904 -46423 955 -46390
rect -9 -46423 42 -46390
rect 655 -46423 706 -46390
rect 489 -46423 540 -46390
rect 904 -46565 955 -46532
rect -9 -46565 42 -46532
rect 655 -46565 706 -46532
rect 489 -46565 540 -46532
rect 738 -46565 789 -46532
rect 904 -46707 955 -46674
rect -9 -46707 42 -46674
rect 406 -46707 457 -46674
rect 904 -46849 955 -46816
rect -9 -46849 42 -46816
rect 406 -46849 457 -46816
rect 738 -46849 789 -46816
rect 904 -46991 955 -46958
rect -9 -46991 42 -46958
rect 406 -46991 457 -46958
rect 655 -46991 706 -46958
rect 904 -47133 955 -47100
rect -9 -47133 42 -47100
rect 655 -47133 706 -47100
rect 406 -47133 457 -47100
rect 738 -47133 789 -47100
rect 904 -47275 955 -47242
rect -9 -47275 42 -47242
rect 406 -47275 457 -47242
rect 489 -47275 540 -47242
rect 904 -47417 955 -47384
rect -9 -47417 42 -47384
rect 406 -47417 457 -47384
rect 489 -47417 540 -47384
rect 738 -47417 789 -47384
rect 904 -47559 955 -47526
rect -9 -47559 42 -47526
rect 406 -47559 457 -47526
rect 655 -47559 706 -47526
rect 489 -47559 540 -47526
rect 904 -47701 955 -47668
rect -9 -47701 42 -47668
rect 655 -47701 706 -47668
rect 489 -47701 540 -47668
rect 406 -47701 457 -47668
rect 738 -47701 789 -47668
rect 904 -47843 955 -47810
rect -9 -47843 42 -47810
rect 240 -47843 291 -47810
rect 904 -47985 955 -47952
rect -9 -47985 42 -47952
rect 240 -47985 291 -47952
rect 738 -47985 789 -47952
rect 904 -48127 955 -48094
rect -9 -48127 42 -48094
rect 655 -48127 706 -48094
rect 240 -48127 291 -48094
rect 904 -48269 955 -48236
rect -9 -48269 42 -48236
rect 655 -48269 706 -48236
rect 240 -48269 291 -48236
rect 738 -48269 789 -48236
rect 904 -48411 955 -48378
rect -9 -48411 42 -48378
rect 489 -48411 540 -48378
rect 240 -48411 291 -48378
rect 904 -48553 955 -48520
rect -9 -48553 42 -48520
rect 489 -48553 540 -48520
rect 240 -48553 291 -48520
rect 738 -48553 789 -48520
rect 904 -48695 955 -48662
rect -9 -48695 42 -48662
rect 655 -48695 706 -48662
rect 489 -48695 540 -48662
rect 240 -48695 291 -48662
rect 904 -48837 955 -48804
rect -9 -48837 42 -48804
rect 655 -48837 706 -48804
rect 489 -48837 540 -48804
rect 240 -48837 291 -48804
rect 738 -48837 789 -48804
rect 904 -48979 955 -48946
rect -9 -48979 42 -48946
rect 406 -48979 457 -48946
rect 240 -48979 291 -48946
rect 904 -49121 955 -49088
rect -9 -49121 42 -49088
rect 406 -49121 457 -49088
rect 240 -49121 291 -49088
rect 738 -49121 789 -49088
rect 904 -49263 955 -49230
rect -9 -49263 42 -49230
rect 406 -49263 457 -49230
rect 655 -49263 706 -49230
rect 240 -49263 291 -49230
rect 904 -49405 955 -49372
rect -9 -49405 42 -49372
rect 655 -49405 706 -49372
rect 406 -49405 457 -49372
rect 240 -49405 291 -49372
rect 738 -49405 789 -49372
rect 904 -49547 955 -49514
rect -9 -49547 42 -49514
rect 406 -49547 457 -49514
rect 489 -49547 540 -49514
rect 240 -49547 291 -49514
rect 904 -49689 955 -49656
rect -9 -49689 42 -49656
rect 406 -49689 457 -49656
rect 489 -49689 540 -49656
rect 240 -49689 291 -49656
rect 738 -49689 789 -49656
rect 904 -49831 955 -49798
rect -9 -49831 42 -49798
rect 406 -49831 457 -49798
rect 655 -49831 706 -49798
rect 489 -49831 540 -49798
rect 240 -49831 291 -49798
rect 904 -49973 955 -49940
rect -9 -49973 42 -49940
rect 655 -49973 706 -49940
rect 489 -49973 540 -49940
rect 406 -49973 457 -49940
rect 240 -49973 291 -49940
rect 738 -49973 789 -49940
rect 904 -50115 955 -50082
rect -9 -50115 42 -50082
rect 157 -50115 208 -50082
rect 904 -50257 955 -50224
rect -9 -50257 42 -50224
rect 157 -50257 208 -50224
rect 738 -50257 789 -50224
rect 904 -50399 955 -50366
rect -9 -50399 42 -50366
rect 655 -50399 706 -50366
rect 157 -50399 208 -50366
rect 904 -50541 955 -50508
rect -9 -50541 42 -50508
rect 655 -50541 706 -50508
rect 157 -50541 208 -50508
rect 738 -50541 789 -50508
rect 904 -50683 955 -50650
rect -9 -50683 42 -50650
rect 489 -50683 540 -50650
rect 157 -50683 208 -50650
rect 904 -50825 955 -50792
rect -9 -50825 42 -50792
rect 489 -50825 540 -50792
rect 157 -50825 208 -50792
rect 738 -50825 789 -50792
rect 904 -50967 955 -50934
rect -9 -50967 42 -50934
rect 655 -50967 706 -50934
rect 489 -50967 540 -50934
rect 157 -50967 208 -50934
rect 904 -51109 955 -51076
rect -9 -51109 42 -51076
rect 655 -51109 706 -51076
rect 489 -51109 540 -51076
rect 157 -51109 208 -51076
rect 738 -51109 789 -51076
rect 904 -51251 955 -51218
rect -9 -51251 42 -51218
rect 406 -51251 457 -51218
rect 157 -51251 208 -51218
rect 904 -51393 955 -51360
rect -9 -51393 42 -51360
rect 406 -51393 457 -51360
rect 157 -51393 208 -51360
rect 738 -51393 789 -51360
rect 904 -51535 955 -51502
rect -9 -51535 42 -51502
rect 406 -51535 457 -51502
rect 655 -51535 706 -51502
rect 157 -51535 208 -51502
rect 904 -51677 955 -51644
rect -9 -51677 42 -51644
rect 655 -51677 706 -51644
rect 406 -51677 457 -51644
rect 157 -51677 208 -51644
rect 738 -51677 789 -51644
rect 904 -51819 955 -51786
rect -9 -51819 42 -51786
rect 406 -51819 457 -51786
rect 489 -51819 540 -51786
rect 157 -51819 208 -51786
rect 904 -51961 955 -51928
rect -9 -51961 42 -51928
rect 406 -51961 457 -51928
rect 489 -51961 540 -51928
rect 157 -51961 208 -51928
rect 738 -51961 789 -51928
rect 904 -52103 955 -52070
rect -9 -52103 42 -52070
rect 406 -52103 457 -52070
rect 655 -52103 706 -52070
rect 489 -52103 540 -52070
rect 157 -52103 208 -52070
rect 904 -52245 955 -52212
rect -9 -52245 42 -52212
rect 655 -52245 706 -52212
rect 489 -52245 540 -52212
rect 406 -52245 457 -52212
rect 157 -52245 208 -52212
rect 738 -52245 789 -52212
rect 904 -52387 955 -52354
rect -9 -52387 42 -52354
rect 240 -52387 291 -52354
rect 157 -52387 208 -52354
rect 904 -52529 955 -52496
rect -9 -52529 42 -52496
rect 240 -52529 291 -52496
rect 157 -52529 208 -52496
rect 738 -52529 789 -52496
rect 904 -52671 955 -52638
rect -9 -52671 42 -52638
rect 655 -52671 706 -52638
rect 240 -52671 291 -52638
rect 157 -52671 208 -52638
rect 904 -52813 955 -52780
rect -9 -52813 42 -52780
rect 655 -52813 706 -52780
rect 240 -52813 291 -52780
rect 157 -52813 208 -52780
rect 738 -52813 789 -52780
rect 904 -52955 955 -52922
rect -9 -52955 42 -52922
rect 489 -52955 540 -52922
rect 240 -52955 291 -52922
rect 157 -52955 208 -52922
rect 904 -53097 955 -53064
rect -9 -53097 42 -53064
rect 489 -53097 540 -53064
rect 240 -53097 291 -53064
rect 157 -53097 208 -53064
rect 738 -53097 789 -53064
rect 904 -53239 955 -53206
rect -9 -53239 42 -53206
rect 655 -53239 706 -53206
rect 489 -53239 540 -53206
rect 240 -53239 291 -53206
rect 157 -53239 208 -53206
rect 904 -53381 955 -53348
rect -9 -53381 42 -53348
rect 655 -53381 706 -53348
rect 489 -53381 540 -53348
rect 240 -53381 291 -53348
rect 157 -53381 208 -53348
rect 738 -53381 789 -53348
rect 904 -53523 955 -53490
rect -9 -53523 42 -53490
rect 406 -53523 457 -53490
rect 240 -53523 291 -53490
rect 157 -53523 208 -53490
rect 904 -53665 955 -53632
rect -9 -53665 42 -53632
rect 406 -53665 457 -53632
rect 240 -53665 291 -53632
rect 157 -53665 208 -53632
rect 738 -53665 789 -53632
rect 904 -53807 955 -53774
rect -9 -53807 42 -53774
rect 406 -53807 457 -53774
rect 655 -53807 706 -53774
rect 240 -53807 291 -53774
rect 157 -53807 208 -53774
rect 904 -53949 955 -53916
rect -9 -53949 42 -53916
rect 655 -53949 706 -53916
rect 406 -53949 457 -53916
rect 240 -53949 291 -53916
rect 157 -53949 208 -53916
rect 738 -53949 789 -53916
rect 904 -54091 955 -54058
rect -9 -54091 42 -54058
rect 406 -54091 457 -54058
rect 489 -54091 540 -54058
rect 240 -54091 291 -54058
rect 157 -54091 208 -54058
rect 904 -54233 955 -54200
rect -9 -54233 42 -54200
rect 406 -54233 457 -54200
rect 489 -54233 540 -54200
rect 240 -54233 291 -54200
rect 157 -54233 208 -54200
rect 738 -54233 789 -54200
rect 904 -54375 955 -54342
rect -9 -54375 42 -54342
rect 406 -54375 457 -54342
rect 655 -54375 706 -54342
rect 489 -54375 540 -54342
rect 240 -54375 291 -54342
rect 157 -54375 208 -54342
rect -9 -54517 42 -54484
rect 655 -54517 706 -54484
rect 489 -54517 540 -54484
rect 406 -54517 457 -54484
rect 240 -54517 291 -54484
rect 157 -54517 208 -54484
rect 738 -54517 789 -54484
rect 904 -54801 955 -54768
rect 904 -54943 955 -54910
rect 738 -55085 789 -55052
rect 904 -55227 955 -55194
rect 655 -55227 706 -55194
rect 738 -55227 789 -55194
rect 904 -55369 955 -55336
rect 655 -55369 706 -55336
rect 904 -55511 955 -55478
rect 655 -55511 706 -55478
rect 738 -55511 789 -55478
rect 904 -55653 955 -55620
rect 489 -55653 540 -55620
rect 738 -55653 789 -55620
rect 904 -55795 955 -55762
rect 655 -55795 706 -55762
rect 489 -55795 540 -55762
rect 738 -55795 789 -55762
rect 904 -55937 955 -55904
rect 655 -55937 706 -55904
rect 489 -55937 540 -55904
rect 738 -55937 789 -55904
rect 904 -56079 955 -56046
rect 406 -56079 457 -56046
rect 738 -56079 789 -56046
rect 904 -56221 955 -56188
rect 406 -56221 457 -56188
rect 655 -56221 706 -56188
rect 904 -56363 955 -56330
rect 655 -56363 706 -56330
rect 406 -56363 457 -56330
rect 489 -56363 540 -56330
rect 738 -56363 789 -56330
rect 904 -56505 955 -56472
rect 406 -56505 457 -56472
rect 489 -56505 540 -56472
rect 655 -56505 706 -56472
rect 738 -56505 789 -56472
rect 904 -56647 955 -56614
rect 655 -56647 706 -56614
rect 489 -56647 540 -56614
rect 406 -56647 457 -56614
rect 240 -56647 291 -56614
rect 738 -56647 789 -56614
rect 904 -56789 955 -56756
rect 655 -56789 706 -56756
rect 240 -56789 291 -56756
rect 738 -56789 789 -56756
rect 489 -56931 540 -56898
rect 240 -56931 291 -56898
rect 738 -56931 789 -56898
rect 904 -57073 955 -57040
rect 655 -57073 706 -57040
rect 489 -57073 540 -57040
rect 240 -57073 291 -57040
rect 738 -57073 789 -57040
rect 904 -57215 955 -57182
rect 406 -57215 457 -57182
rect 655 -57215 706 -57182
rect 240 -57215 291 -57182
rect 904 -57357 955 -57324
rect 655 -57357 706 -57324
rect 406 -57357 457 -57324
rect 240 -57357 291 -57324
rect 489 -57357 540 -57324
rect 738 -57357 789 -57324
rect 904 -57499 955 -57466
rect 406 -57499 457 -57466
rect 489 -57499 540 -57466
rect 655 -57499 706 -57466
rect 240 -57499 291 -57466
rect 738 -57499 789 -57466
rect 904 -57641 955 -57608
rect 157 -57641 208 -57608
rect 738 -57641 789 -57608
rect 904 -57783 955 -57750
rect 655 -57783 706 -57750
rect 489 -57783 540 -57750
rect 157 -57783 208 -57750
rect 738 -57783 789 -57750
rect 904 -57925 955 -57892
rect 655 -57925 706 -57892
rect 489 -57925 540 -57892
rect 157 -57925 208 -57892
rect 738 -57925 789 -57892
rect 904 -58067 955 -58034
rect 406 -58067 457 -58034
rect 655 -58067 706 -58034
rect 157 -58067 208 -58034
rect 738 -58067 789 -58034
rect 406 -58209 457 -58176
rect 489 -58209 540 -58176
rect 157 -58209 208 -58176
rect 738 -58209 789 -58176
rect 904 -58351 955 -58318
rect 655 -58351 706 -58318
rect 489 -58351 540 -58318
rect 406 -58351 457 -58318
rect 240 -58351 291 -58318
rect 157 -58351 208 -58318
rect 904 -58493 955 -58460
rect 655 -58493 706 -58460
rect 240 -58493 291 -58460
rect 157 -58493 208 -58460
rect 738 -58493 789 -58460
rect 904 -58635 955 -58602
rect 489 -58635 540 -58602
rect 655 -58635 706 -58602
rect 240 -58635 291 -58602
rect 157 -58635 208 -58602
rect 738 -58635 789 -58602
rect 904 -58777 955 -58744
rect 406 -58777 457 -58744
rect 240 -58777 291 -58744
rect 157 -58777 208 -58744
rect 738 -58777 789 -58744
rect 904 -58919 955 -58886
rect 489 -58919 540 -58886
rect 655 -58919 706 -58886
rect 406 -58919 457 -58886
rect 240 -58919 291 -58886
rect 157 -58919 208 -58886
rect 738 -58919 789 -58886
rect -9 -59061 42 -59028
rect 406 -59061 457 -59028
rect 655 -59061 706 -59028
rect 489 -59061 540 -59028
rect 240 -59061 291 -59028
rect 157 -59061 208 -59028
rect 904 -59203 955 -59170
rect -9 -59203 42 -59170
rect 655 -59203 706 -59170
rect 738 -59203 789 -59170
rect 904 -59345 955 -59312
rect -9 -59345 42 -59312
rect 655 -59345 706 -59312
rect 489 -59345 540 -59312
rect 904 -59487 955 -59454
rect -9 -59487 42 -59454
rect 655 -59487 706 -59454
rect 489 -59487 540 -59454
rect 406 -59487 457 -59454
rect 738 -59487 789 -59454
rect 904 -59629 955 -59596
rect -9 -59629 42 -59596
rect 406 -59629 457 -59596
rect 655 -59629 706 -59596
rect 489 -59629 540 -59596
rect 904 -59771 955 -59738
rect -9 -59771 42 -59738
rect 406 -59771 457 -59738
rect 489 -59771 540 -59738
rect 655 -59771 706 -59738
rect 738 -59771 789 -59738
rect 904 -59913 955 -59880
rect -9 -59913 42 -59880
rect 655 -59913 706 -59880
rect 240 -59913 291 -59880
rect 738 -59913 789 -59880
rect 904 -60055 955 -60022
rect -9 -60055 42 -60022
rect 655 -60055 706 -60022
rect 489 -60055 540 -60022
rect 240 -60055 291 -60022
rect 738 -60055 789 -60022
rect 904 -60197 955 -60164
rect -9 -60197 42 -60164
rect 655 -60197 706 -60164
rect 489 -60197 540 -60164
rect 406 -60197 457 -60164
rect 240 -60197 291 -60164
rect 904 -60339 955 -60306
rect -9 -60339 42 -60306
rect 406 -60339 457 -60306
rect 655 -60339 706 -60306
rect 240 -60339 291 -60306
rect 738 -60339 789 -60306
rect 904 -60481 955 -60448
rect -9 -60481 42 -60448
rect 406 -60481 457 -60448
rect 489 -60481 540 -60448
rect 655 -60481 706 -60448
rect 240 -60481 291 -60448
rect 904 -60623 955 -60590
rect -9 -60623 42 -60590
rect 655 -60623 706 -60590
rect 489 -60623 540 -60590
rect 406 -60623 457 -60590
rect 240 -60623 291 -60590
rect 157 -60623 208 -60590
rect 738 -60623 789 -60590
rect -9 -60765 42 -60732
rect 655 -60765 706 -60732
rect 157 -60765 208 -60732
rect 738 -60765 789 -60732
rect 904 -60907 955 -60874
rect -9 -60907 42 -60874
rect 489 -60907 540 -60874
rect 157 -60907 208 -60874
rect 738 -60907 789 -60874
rect -9 -61049 42 -61016
rect 655 -61049 706 -61016
rect 489 -61049 540 -61016
rect 406 -61049 457 -61016
rect 157 -61049 208 -61016
rect 738 -61049 789 -61016
rect 904 -61191 955 -61158
rect -9 -61191 42 -61158
rect 406 -61191 457 -61158
rect 655 -61191 706 -61158
rect 157 -61191 208 -61158
rect 738 -61191 789 -61158
rect 904 -61333 955 -61300
rect -9 -61333 42 -61300
rect 655 -61333 706 -61300
rect 406 -61333 457 -61300
rect 157 -61333 208 -61300
rect 738 -61333 789 -61300
rect 489 -61333 540 -61300
rect -9 -61475 42 -61442
rect 406 -61475 457 -61442
rect 655 -61475 706 -61442
rect 489 -61475 540 -61442
rect 157 -61475 208 -61442
rect 738 -61475 789 -61442
rect -9 -61617 42 -61584
rect 240 -61617 291 -61584
rect 157 -61617 208 -61584
rect 738 -61617 789 -61584
rect -9 -61759 42 -61726
rect 655 -61759 706 -61726
rect 240 -61759 291 -61726
rect 157 -61759 208 -61726
rect 738 -61759 789 -61726
rect -9 -61901 42 -61868
rect 489 -61901 540 -61868
rect 240 -61901 291 -61868
rect 157 -61901 208 -61868
rect 738 -61901 789 -61868
rect 904 -62043 955 -62010
rect -9 -62043 42 -62010
rect 489 -62043 540 -62010
rect 655 -62043 706 -62010
rect 240 -62043 291 -62010
rect 157 -62043 208 -62010
rect 738 -62043 789 -62010
rect -9 -62185 42 -62152
rect 655 -62185 706 -62152
rect 489 -62185 540 -62152
rect 240 -62185 291 -62152
rect 157 -62185 208 -62152
rect 738 -62185 789 -62152
rect 406 -62185 457 -62152
rect 904 -62327 955 -62294
rect -9 -62327 42 -62294
rect 406 -62327 457 -62294
rect 240 -62327 291 -62294
rect 157 -62327 208 -62294
rect 738 -62327 789 -62294
rect 904 -62469 955 -62436
rect -9 -62469 42 -62436
rect 406 -62469 457 -62436
rect 655 -62469 706 -62436
rect 240 -62469 291 -62436
rect 157 -62469 208 -62436
rect -9 -62611 42 -62578
rect 655 -62611 706 -62578
rect 406 -62611 457 -62578
rect 240 -62611 291 -62578
rect 157 -62611 208 -62578
rect 738 -62611 789 -62578
rect 489 -62611 540 -62578
rect 904 -62753 955 -62720
rect -9 -62753 42 -62720
rect 406 -62753 457 -62720
rect 489 -62753 540 -62720
rect 240 -62753 291 -62720
rect 157 -62753 208 -62720
rect 738 -62753 789 -62720
rect 904 -62895 955 -62862
rect -9 -62895 42 -62862
rect 406 -62895 457 -62862
rect 489 -62895 540 -62862
rect 240 -62895 291 -62862
rect 157 -62895 208 -62862
rect 738 -62895 789 -62862
rect 904 -63037 955 -63004
rect -9 -63037 42 -63004
rect 406 -63037 457 -63004
rect 655 -63037 706 -63004
rect 489 -63037 540 -63004
rect 240 -63037 291 -63004
rect 157 -63037 208 -63004
rect 904 -63179 955 -63146
rect -9 -63179 42 -63146
rect 655 -63179 706 -63146
rect 489 -63179 540 -63146
rect 406 -63179 457 -63146
rect 240 -63179 291 -63146
rect 157 -63179 208 -63146
rect 738 -63179 789 -63146
rect -9 -63321 42 -63288
rect 655 -63321 706 -63288
rect 489 -63321 540 -63288
rect 406 -63321 457 -63288
rect 240 -63321 291 -63288
rect 157 -63321 208 -63288
rect 738 -63321 789 -63288
rect 904 -63463 955 -63430
rect -9 -63463 42 -63430
rect 655 -63463 706 -63430
rect 489 -63463 540 -63430
rect 406 -63463 457 -63430
rect 240 -63463 291 -63430
rect 157 -63463 208 -63430
rect 738 -63463 789 -63430
rect 904 -63605 955 -63572
rect -9 -63605 42 -63572
rect 655 -63605 706 -63572
rect 489 -63605 540 -63572
rect 406 -63605 457 -63572
rect 240 -63605 291 -63572
rect 157 -63605 208 -63572
rect 738 -63605 789 -63572
rect 904 -63747 955 -63714
rect -9 -63747 42 -63714
rect 655 -63747 706 -63714
rect 489 -63747 540 -63714
rect 406 -63747 457 -63714
rect 240 -63747 291 -63714
rect 157 -63747 208 -63714
rect 738 -63747 789 -63714
rect 904 -63889 955 -63856
rect -9 -63889 42 -63856
rect 655 -63889 706 -63856
rect 489 -63889 540 -63856
rect 406 -63889 457 -63856
rect 240 -63889 291 -63856
rect 157 -63889 208 -63856
rect 738 -63889 789 -63856
rect -9 -64031 42 -63998
rect 655 -64031 706 -63998
rect 489 -64031 540 -63998
rect 406 -64031 457 -63998
rect 240 -64031 291 -63998
rect 157 -64031 208 -63998
rect 738 -64031 789 -63998
rect 904 -64173 955 -64140
rect -9 -64173 42 -64140
rect 655 -64173 706 -64140
rect 489 -64173 540 -64140
rect 406 -64173 457 -64140
rect 240 -64173 291 -64140
rect 157 -64173 208 -64140
rect 904 -64315 955 -64282
rect -9 -64315 42 -64282
rect 406 -64315 457 -64282
rect 655 -64315 706 -64282
rect 489 -64315 540 -64282
rect 240 -64315 291 -64282
rect 157 -64315 208 -64282
rect 738 -64315 789 -64282
rect -9 -64457 42 -64424
rect 406 -64457 457 -64424
rect 489 -64457 540 -64424
rect 240 -64457 291 -64424
rect 157 -64457 208 -64424
rect 738 -64457 789 -64424
rect 904 -64599 955 -64566
rect -9 -64599 42 -64566
rect 406 -64599 457 -64566
rect 489 -64599 540 -64566
rect 240 -64599 291 -64566
rect 157 -64599 208 -64566
rect 904 -64741 955 -64708
rect -9 -64741 42 -64708
rect 655 -64741 706 -64708
rect 406 -64741 457 -64708
rect 240 -64741 291 -64708
rect 157 -64741 208 -64708
rect 738 -64741 789 -64708
rect 904 -64883 955 -64850
rect -9 -64883 42 -64850
rect 406 -64883 457 -64850
rect 655 -64883 706 -64850
rect 240 -64883 291 -64850
rect 157 -64883 208 -64850
rect 738 -64883 789 -64850
rect 904 -65025 955 -64992
rect -9 -65025 42 -64992
rect 406 -65025 457 -64992
rect 240 -65025 291 -64992
rect 157 -65025 208 -64992
rect 904 -65167 955 -65134
rect -9 -65167 42 -65134
rect 655 -65167 706 -65134
rect 489 -65167 540 -65134
rect 240 -65167 291 -65134
rect 157 -65167 208 -65134
rect 738 -65167 789 -65134
rect 904 -65309 955 -65276
rect -9 -65309 42 -65276
rect 489 -65309 540 -65276
rect 240 -65309 291 -65276
rect 157 -65309 208 -65276
rect 738 -65309 789 -65276
rect -9 -65451 42 -65418
rect 489 -65451 540 -65418
rect 655 -65451 706 -65418
rect 240 -65451 291 -65418
rect 157 -65451 208 -65418
rect 738 -65451 789 -65418
rect -9 -65593 42 -65560
rect 655 -65593 706 -65560
rect 240 -65593 291 -65560
rect 157 -65593 208 -65560
rect 738 -65593 789 -65560
rect -9 -65735 42 -65702
rect 655 -65735 706 -65702
rect 489 -65735 540 -65702
rect 240 -65735 291 -65702
rect 157 -65735 208 -65702
rect 738 -65735 789 -65702
rect 406 -65735 457 -65702
rect -9 -65877 42 -65844
rect 406 -65877 457 -65844
rect 655 -65877 706 -65844
rect 489 -65877 540 -65844
rect 157 -65877 208 -65844
rect 738 -65877 789 -65844
rect 904 -66019 955 -65986
rect -9 -66019 42 -65986
rect 655 -66019 706 -65986
rect 406 -66019 457 -65986
rect 157 -66019 208 -65986
rect 738 -66019 789 -65986
rect 904 -66161 955 -66128
rect -9 -66161 42 -66128
rect 406 -66161 457 -66128
rect 157 -66161 208 -66128
rect 738 -66161 789 -66128
rect 904 -66303 955 -66270
rect -9 -66303 42 -66270
rect 655 -66303 706 -66270
rect 489 -66303 540 -66270
rect 157 -66303 208 -66270
rect 738 -66303 789 -66270
rect 904 -66445 955 -66412
rect -9 -66445 42 -66412
rect 489 -66445 540 -66412
rect 655 -66445 706 -66412
rect 157 -66445 208 -66412
rect 738 -66445 789 -66412
rect 904 -66587 955 -66554
rect -9 -66587 42 -66554
rect 655 -66587 706 -66554
rect 157 -66587 208 -66554
rect -9 -66729 42 -66696
rect 655 -66729 706 -66696
rect 489 -66729 540 -66696
rect 406 -66729 457 -66696
rect 240 -66729 291 -66696
rect 738 -66729 789 -66696
rect 904 -66871 955 -66838
rect -9 -66871 42 -66838
rect 406 -66871 457 -66838
rect 489 -66871 540 -66838
rect 655 -66871 706 -66838
rect 240 -66871 291 -66838
rect 738 -66871 789 -66838
rect 904 -67013 955 -66980
rect -9 -67013 42 -66980
rect 406 -67013 457 -66980
rect 240 -67013 291 -66980
rect 738 -67013 789 -66980
rect 904 -67155 955 -67122
rect -9 -67155 42 -67122
rect 655 -67155 706 -67122
rect 489 -67155 540 -67122
rect 240 -67155 291 -67122
rect 738 -67155 789 -67122
rect 904 -67297 955 -67264
rect -9 -67297 42 -67264
rect 655 -67297 706 -67264
rect 240 -67297 291 -67264
rect 738 -67297 789 -67264
rect -9 -67439 42 -67406
rect 655 -67439 706 -67406
rect 489 -67439 540 -67406
rect 406 -67439 457 -67406
rect 240 -67439 291 -67406
rect 738 -67439 789 -67406
rect 904 -67581 955 -67548
rect -9 -67581 42 -67548
rect 406 -67581 457 -67548
rect 489 -67581 540 -67548
rect 738 -67581 789 -67548
rect 904 -67723 955 -67690
rect -9 -67723 42 -67690
rect 406 -67723 457 -67690
rect 655 -67723 706 -67690
rect 738 -67723 789 -67690
rect 904 -67865 955 -67832
rect -9 -67865 42 -67832
rect 655 -67865 706 -67832
rect 489 -67865 540 -67832
rect 738 -67865 789 -67832
rect 904 -68007 955 -67974
rect -9 -68007 42 -67974
rect 655 -68007 706 -67974
rect 489 -68007 540 -67974
rect 738 -68007 789 -67974
rect 904 -68149 955 -68116
rect -9 -68149 42 -68116
rect 738 -68149 789 -68116
rect 904 -68291 955 -68258
rect 406 -68291 457 -68258
rect 655 -68291 706 -68258
rect 489 -68291 540 -68258
rect 240 -68291 291 -68258
rect 157 -68291 208 -68258
rect 904 -68433 955 -68400
rect 655 -68433 706 -68400
rect 406 -68433 457 -68400
rect 240 -68433 291 -68400
rect 157 -68433 208 -68400
rect 738 -68433 789 -68400
rect 904 -68575 955 -68542
rect 406 -68575 457 -68542
rect 655 -68575 706 -68542
rect 489 -68575 540 -68542
rect 240 -68575 291 -68542
rect 157 -68575 208 -68542
rect 904 -68717 955 -68684
rect 489 -68717 540 -68684
rect 655 -68717 706 -68684
rect 240 -68717 291 -68684
rect 157 -68717 208 -68684
rect 738 -68717 789 -68684
rect 904 -68859 955 -68826
rect 655 -68859 706 -68826
rect 240 -68859 291 -68826
rect 157 -68859 208 -68826
rect 904 -69001 955 -68968
rect 655 -69001 706 -68968
rect 489 -69001 540 -68968
rect 406 -69001 457 -68968
rect 157 -69001 208 -68968
rect 738 -69001 789 -68968
rect 904 -69143 955 -69110
rect 406 -69143 457 -69110
rect 489 -69143 540 -69110
rect 655 -69143 706 -69110
rect 157 -69143 208 -69110
rect 904 -69285 955 -69252
rect 406 -69285 457 -69252
rect 655 -69285 706 -69252
rect 489 -69285 540 -69252
rect 157 -69285 208 -69252
rect 738 -69285 789 -69252
rect 904 -69427 955 -69394
rect 655 -69427 706 -69394
rect 489 -69427 540 -69394
rect 157 -69427 208 -69394
rect 904 -69569 955 -69536
rect 655 -69569 706 -69536
rect 157 -69569 208 -69536
rect 738 -69569 789 -69536
rect 904 -69711 955 -69678
rect 240 -69711 291 -69678
rect 655 -69711 706 -69678
rect 489 -69711 540 -69678
rect 406 -69711 457 -69678
rect 157 -69711 208 -69678
rect 738 -69711 789 -69678
rect 904 -69853 955 -69820
rect 406 -69853 457 -69820
rect 489 -69853 540 -69820
rect 240 -69853 291 -69820
rect 738 -69853 789 -69820
rect 655 -69995 706 -69962
rect 406 -69995 457 -69962
rect 240 -69995 291 -69962
rect 738 -69995 789 -69962
rect 904 -70137 955 -70104
rect 406 -70137 457 -70104
rect 655 -70137 706 -70104
rect 240 -70137 291 -70104
rect 489 -70137 540 -70104
rect 738 -70137 789 -70104
rect 655 -70279 706 -70246
rect 489 -70279 540 -70246
rect 240 -70279 291 -70246
rect 738 -70279 789 -70246
rect 904 -70421 955 -70388
rect 655 -70421 706 -70388
rect 489 -70421 540 -70388
rect 240 -70421 291 -70388
rect 904 -70563 955 -70530
rect 240 -70563 291 -70530
rect 738 -70563 789 -70530
rect 904 -70705 955 -70672
rect 655 -70705 706 -70672
rect 489 -70705 540 -70672
rect 406 -70705 457 -70672
rect 738 -70705 789 -70672
rect 904 -70847 955 -70814
rect 406 -70847 457 -70814
rect 489 -70847 540 -70814
rect 738 -70847 789 -70814
rect 904 -70989 955 -70956
rect 655 -70989 706 -70956
rect 406 -70989 457 -70956
rect 738 -70989 789 -70956
rect 406 -71131 457 -71098
rect 655 -71131 706 -71098
rect 738 -71131 789 -71098
rect 904 -71273 955 -71240
rect 406 -71273 457 -71240
rect 655 -71273 706 -71240
rect 489 -71273 540 -71240
rect 738 -71273 789 -71240
rect 655 -71415 706 -71382
rect 489 -71415 540 -71382
rect 738 -71415 789 -71382
rect 904 -71557 955 -71524
rect 489 -71557 540 -71524
rect 738 -71557 789 -71524
rect 904 -71699 955 -71666
rect 655 -71699 706 -71666
rect 489 -71699 540 -71666
rect 738 -71699 789 -71666
rect 904 -71841 955 -71808
rect 655 -71841 706 -71808
rect 738 -71841 789 -71808
rect 904 -71983 955 -71950
rect 655 -71983 706 -71950
rect 738 -72125 789 -72092
rect 904 -72125 955 -72092
rect 904 -72267 955 -72234
rect 738 -72267 789 -72234
rect 904 -72409 955 -72376
rect 904 -36095 955 -36057
rect 904 -29208 955 -29170
rect 904 -29634 955 -29596
rect 904 -10535 955 -10497
rect 904 -42911 955 -42873
rect 904 -66980 955 -66942
rect 904 -42627 955 -42589
rect 904 -15363 955 -15325
rect 904 -26013 955 -25975
rect 904 -34675 955 -34637
rect 904 -41633 955 -41595
rect 904 -20901 955 -20863
rect 904 -30628 955 -30590
rect 904 -57182 955 -57144
rect 904 -43053 955 -43015
rect 904 -11245 955 -11207
rect 904 -41349 955 -41311
rect 904 -71950 955 -71912
rect 904 -28143 955 -28105
rect 904 -31338 955 -31300
rect 904 -56827 955 -56789
rect 904 -37941 955 -37903
rect 904 -31977 955 -31939
rect 904 -68116 955 -68078
rect 904 -27788 955 -27750
rect 904 -15008 955 -14970
rect 904 -70743 955 -70705
rect 904 -16144 955 -16106
rect 904 -10819 955 -10781
rect 904 -59951 955 -59913
rect 904 -43195 955 -43157
rect 904 -24806 955 -24768
rect 904 -22463 955 -22425
rect 904 -9257 955 -9219
rect 904 -62933 955 -62895
rect 904 -58957 955 -58919
rect 904 -13304 955 -13266
rect 904 -33184 955 -33146
rect 904 -20688 955 -20650
rect 904 -67974 955 -67936
rect 904 -24451 955 -24413
rect 904 -49727 955 -49689
rect 904 -10180 955 -10142
rect 904 -57395 955 -57357
rect 904 -29350 955 -29312
rect 904 -23457 955 -23419
rect 904 -25374 955 -25336
rect 904 -11742 955 -11704
rect 904 -35527 955 -35489
rect 904 -16357 955 -16319
rect 904 -24025 955 -23987
rect 904 -25729 955 -25691
rect 904 -20759 955 -20721
rect 904 -35953 955 -35915
rect 904 -66341 955 -66303
rect 904 -13517 955 -13479
rect 904 -53845 955 -53807
rect 904 -62365 955 -62327
rect 904 -17280 955 -17242
rect 904 -49585 955 -49547
rect 904 -43479 955 -43441
rect 904 -31551 955 -31513
rect 904 -22037 955 -21999
rect 904 -27291 955 -27253
rect 904 -65986 955 -65948
rect 904 -47313 955 -47275
rect 904 -35740 955 -35702
rect 904 -38935 955 -38897
rect 904 -28072 955 -28034
rect 904 -55336 955 -55298
rect 904 -20333 955 -20295
rect 904 -51005 955 -50967
rect 904 -15718 955 -15680
rect 904 -52567 955 -52529
rect 904 -19055 955 -19017
rect 904 -30060 955 -30022
rect 904 -54271 955 -54233
rect 904 -35172 955 -35134
rect 904 -50579 955 -50541
rect 904 -31693 955 -31655
rect 904 -43905 955 -43867
rect 904 -70885 955 -70847
rect 904 -12594 955 -12556
rect 904 -26297 955 -26259
rect 904 -62507 955 -62469
rect 904 -19694 955 -19656
rect 904 -64353 955 -64315
rect 904 -14440 955 -14402
rect 904 -46035 955 -45997
rect 904 -24877 955 -24839
rect 904 -27930 955 -27892
rect 904 -28853 955 -28815
rect 904 -35385 955 -35347
rect 904 -9683 955 -9645
rect 904 -56330 955 -56292
rect 904 -70956 955 -70918
rect 904 -10464 955 -10426
rect 904 -20546 955 -20508
rect 904 -50863 955 -50825
rect 904 -59738 955 -59700
rect 904 -59170 955 -59132
rect 904 -60874 955 -60836
rect 904 -15292 955 -15254
rect 904 -46461 955 -46423
rect 904 -38651 955 -38613
rect 904 -56046 955 -56008
rect 904 -41065 955 -41027
rect 904 -12736 955 -12698
rect 904 -46177 955 -46139
rect 904 -25516 955 -25478
rect 904 -34746 955 -34708
rect 904 -36166 955 -36128
rect 904 -35314 955 -35276
rect 904 -26510 955 -26472
rect 904 -30841 955 -30803
rect 904 -34959 955 -34921
rect 904 -54981 955 -54943
rect 904 -33397 955 -33359
rect 904 -47455 955 -47417
rect 904 -52283 955 -52245
rect 904 -29563 955 -29525
rect 904 -48733 955 -48695
rect 904 -44615 955 -44577
rect 904 -32971 955 -32933
rect 904 -40355 955 -40317
rect 904 -27646 955 -27608
rect 904 -15576 955 -15538
rect 904 -41917 955 -41879
rect 904 -68755 955 -68717
rect 904 -29776 955 -29738
rect 904 -32758 955 -32720
rect 904 -39645 955 -39607
rect 904 -50721 955 -50683
rect 904 -32687 955 -32649
rect 904 -21753 955 -21715
rect 904 -31764 955 -31726
rect 904 -17564 955 -17526
rect 904 -55762 955 -55724
rect 904 -65276 955 -65238
rect 904 -11032 955 -10994
rect 904 -63146 955 -63108
rect 904 -50153 955 -50115
rect 904 -58531 955 -58493
rect 904 -30912 955 -30874
rect 904 -14511 955 -14473
rect 904 -22605 955 -22567
rect 904 -21966 955 -21928
rect 904 -68471 955 -68433
rect 904 -68968 955 -68930
rect 904 -17990 955 -17952
rect 904 -27504 955 -27466
rect 904 -29989 955 -29951
rect 904 -54839 955 -54801
rect 904 -32474 955 -32436
rect 904 -62720 955 -62682
rect 904 -35598 955 -35560
rect 904 -63856 955 -63818
rect 904 -11103 955 -11065
rect 904 -35882 955 -35844
rect 904 -14866 955 -14828
rect 904 -21469 955 -21431
rect 904 -23599 955 -23561
rect 904 -62081 955 -62043
rect 904 -11884 955 -11846
rect 904 -49017 955 -48979
rect 904 -55549 955 -55511
rect 904 -55620 955 -55582
rect 904 -11529 955 -11491
rect 904 -15434 955 -15396
rect 904 -32403 955 -32365
rect 904 -17209 955 -17171
rect 904 -47881 955 -47843
rect 904 -48449 955 -48411
rect 904 -51715 955 -51677
rect 904 -33894 955 -33856
rect 904 -18771 955 -18733
rect 904 -25587 955 -25549
rect 904 -68613 955 -68575
rect 904 -44473 955 -44435
rect 904 -72092 955 -72054
rect 904 -9825 955 -9787
rect 904 -52141 955 -52103
rect 904 -70459 955 -70421
rect 904 -19126 955 -19088
rect 904 -12807 955 -12769
rect 904 -21185 955 -21147
rect 904 -32261 955 -32223
rect 904 -44189 955 -44151
rect 904 -33539 955 -33501
rect 904 -25019 955 -24981
rect 904 -40781 955 -40743
rect 904 -63643 955 -63605
rect 904 -25232 955 -25194
rect 904 -39077 955 -39039
rect 904 -56543 955 -56505
rect 904 -19907 955 -19869
rect 904 -26936 955 -26898
rect 904 -57466 955 -57428
rect 904 -18629 955 -18591
rect 904 -33681 955 -33643
rect 904 -10677 955 -10639
rect 904 -65205 955 -65167
rect 904 -13588 955 -13550
rect 904 -22747 955 -22709
rect 904 -32190 955 -32152
rect 904 -29847 955 -29809
rect 904 -48023 955 -47985
rect 904 -27717 955 -27679
rect 904 -50437 955 -50399
rect 904 -62010 955 -61972
rect 904 -71879 955 -71841
rect 904 -44899 955 -44861
rect 904 -21398 955 -21360
rect 904 -22818 955 -22780
rect 904 -58389 955 -58351
rect 904 -40497 955 -40459
rect 904 -17422 955 -17384
rect 904 -24096 955 -24058
rect 904 -30131 955 -30093
rect 904 -22534 955 -22496
rect 904 -45183 955 -45145
rect 904 -45467 955 -45429
rect 904 -60164 955 -60126
rect 904 -28640 955 -28602
rect 904 -23741 955 -23703
rect 904 -60306 955 -60268
rect 904 -24593 955 -24555
rect 904 -29066 955 -29028
rect 904 -23173 955 -23135
rect 904 -14937 955 -14899
rect 904 -32545 955 -32507
rect 904 -20475 955 -20437
rect 904 -21682 955 -21644
rect 904 -10890 955 -10852
rect 904 -18132 955 -18094
rect 904 -14724 955 -14686
rect 904 -49301 955 -49263
rect 904 -10748 955 -10710
rect 904 -33610 955 -33572
rect 904 -12239 955 -12201
rect 904 -33965 955 -33927
rect 904 -24380 955 -24342
rect 904 -37231 955 -37193
rect 904 -41775 955 -41737
rect 904 -42201 955 -42163
rect 904 -19268 955 -19230
rect 904 -33823 955 -33785
rect 904 -19410 955 -19372
rect 904 -39929 955 -39891
rect 904 -45609 955 -45571
rect 904 -41491 955 -41453
rect 904 -18416 955 -18378
rect 904 -25090 955 -25052
rect 904 -22179 955 -22141
rect 904 -69891 955 -69853
rect 904 -24735 955 -24697
rect 904 -39503 955 -39465
rect 904 -19481 955 -19443
rect 904 -40071 955 -40033
rect 904 -26652 955 -26614
rect 904 -23244 955 -23206
rect 904 -21043 955 -21005
rect 904 -56685 955 -56647
rect 904 -10393 955 -10355
rect 904 -26368 955 -26330
rect 904 -29705 955 -29667
rect 904 -31835 955 -31797
rect 904 -51289 955 -51251
rect 904 -29279 955 -29241
rect 904 -9470 955 -9432
rect 904 -11671 955 -11633
rect 904 -48165 955 -48127
rect 904 -19197 955 -19159
rect 904 -13943 955 -13905
rect 904 -53419 955 -53381
rect 904 -30770 955 -30732
rect 904 -14298 955 -14260
rect 904 -23315 955 -23277
rect 904 -32048 955 -32010
rect 904 -35669 955 -35631
rect 904 -31622 955 -31584
rect 904 -27078 955 -27040
rect 904 -25871 955 -25833
rect 904 -24167 955 -24129
rect 904 -29137 955 -29099
rect 904 -45751 955 -45713
rect 904 -11955 955 -11917
rect 904 -37515 955 -37477
rect 904 -59596 955 -59558
rect 904 -14014 955 -13976
rect 904 -22676 955 -22638
rect 904 -38509 955 -38471
rect 904 -17848 955 -17810
rect 904 -54910 955 -54872
rect 904 -35030 955 -34992
rect 904 -60022 955 -59984
rect 904 -14369 955 -14331
rect 904 -34249 955 -34211
rect 904 -24309 955 -24271
rect 904 -47171 955 -47133
rect 904 -28427 955 -28389
rect 904 -15150 955 -15112
rect 904 -15221 955 -15183
rect 904 -59312 955 -59274
rect 904 -25800 955 -25762
rect 904 -70530 955 -70492
rect 904 -56401 955 -56363
rect 904 -57608 955 -57570
rect 904 -36947 955 -36909
rect 904 -16712 955 -16674
rect 904 -58318 955 -58280
rect 904 -50295 955 -50257
rect 904 -9328 955 -9290
rect 904 -12026 955 -11988
rect 904 -21114 955 -21076
rect 904 -18984 955 -18946
rect 904 -33042 955 -33004
rect 904 -9541 955 -9503
rect 904 -11387 955 -11349
rect 904 -71311 955 -71273
rect 904 -31196 955 -31158
rect 904 -64566 955 -64528
rect 904 -14227 955 -14189
rect 904 -24238 955 -24200
rect 904 -26581 955 -26543
rect 904 -15505 955 -15467
rect 904 -45041 955 -45003
rect 904 -18558 955 -18520
rect 904 -16286 955 -16248
rect 904 -32332 955 -32294
rect 904 -22889 955 -22851
rect 904 -60661 955 -60623
rect 904 -26723 955 -26685
rect 904 -63501 955 -63463
rect 904 -16925 955 -16887
rect 904 -48591 955 -48553
rect 904 -37799 955 -37761
rect 904 -41207 955 -41169
rect 904 -71666 955 -71628
rect 904 -68897 955 -68859
rect 904 -40639 955 -40601
rect 904 -10251 955 -10213
rect 904 -60945 955 -60907
rect 904 -67548 955 -67510
rect 904 -40213 955 -40175
rect 904 -34178 955 -34140
rect 904 -12878 955 -12840
rect 904 -36663 955 -36625
rect 904 -70672 955 -70634
rect 904 -63714 955 -63676
rect 904 -18061 955 -18023
rect 904 -9754 955 -9716
rect 904 -21824 955 -21786
rect 904 -30699 955 -30661
rect 904 -45893 955 -45855
rect 904 -61158 955 -61120
rect 904 -25942 955 -25904
rect 904 -53703 955 -53665
rect 904 -40923 955 -40885
rect 904 -56614 955 -56576
rect 904 -16428 955 -16390
rect 904 -35101 955 -35063
rect 904 -50011 955 -49973
rect 904 -10109 955 -10071
rect 904 -13233 955 -13195
rect 904 -12452 955 -12414
rect 904 -34604 955 -34566
rect 904 -13446 955 -13408
rect 904 -57679 955 -57641
rect 904 -13375 955 -13337
rect 904 -34320 955 -34282
rect 904 -16641 955 -16603
rect 904 -16570 955 -16532
rect 904 -31409 955 -31371
rect 904 -17493 955 -17455
rect 904 -64779 955 -64741
rect 904 -23102 955 -23064
rect 904 -53561 955 -53523
rect 904 -27575 955 -27537
rect 904 -29421 955 -29383
rect 904 -62294 955 -62256
rect 904 -46887 955 -46849
rect 904 -53987 955 -53949
rect 904 -57963 955 -57925
rect 904 -36024 955 -35986
rect 904 -32900 955 -32862
rect 904 -30486 955 -30448
rect 904 -45325 955 -45287
rect 904 -33468 955 -33430
rect 904 -22321 955 -22283
rect 904 -15789 955 -15751
rect 904 -17067 955 -17029
rect 904 -28995 955 -28957
rect 904 -52851 955 -52813
rect 904 -23670 955 -23632
rect 904 -30344 955 -30306
rect 904 -69323 955 -69285
rect 904 -20404 955 -20366
rect 904 -24948 955 -24910
rect 904 -26155 955 -26117
rect 904 -31125 955 -31087
rect 904 -28214 955 -28176
rect 904 -32616 955 -32578
rect 904 -27859 955 -27821
rect 904 -15079 955 -15041
rect 904 -70814 955 -70776
rect 904 -25303 955 -25265
rect 904 -13730 955 -13692
rect 904 -23031 955 -22993
rect 904 -70601 955 -70563
rect 904 -27362 955 -27324
rect 904 -39361 955 -39323
rect 904 -16215 955 -16177
rect 904 -25445 955 -25407
rect 904 -37089 955 -37051
rect 904 -57821 955 -57783
rect 904 -19552 955 -19514
rect 904 -28782 955 -28744
rect 904 -39219 955 -39181
rect 904 -19623 955 -19585
rect 904 -70104 955 -70066
rect 904 -66128 955 -66090
rect 904 -51857 955 -51819
rect 904 -56472 955 -56434
rect 904 -63430 955 -63392
rect 904 -16073 955 -16035
rect 904 -10322 955 -10284
rect 904 -64921 955 -64883
rect 904 -58815 955 -58777
rect 904 -18700 955 -18662
rect 904 -28498 955 -28460
rect 904 -71524 955 -71486
rect 904 -36308 955 -36270
rect 904 -31054 955 -31016
rect 904 -67335 955 -67297
rect 904 -57111 955 -57073
rect 904 -26226 955 -26188
rect 904 -61229 955 -61191
rect 904 -67690 955 -67652
rect 904 -21895 955 -21857
rect 904 -9612 955 -9574
rect 904 -69181 955 -69143
rect 904 -67122 955 -67084
rect 904 -67832 955 -67794
rect 904 -24522 955 -24484
rect 904 -63785 955 -63747
rect 904 -30983 955 -30945
rect 904 -17777 955 -17739
rect 904 -52425 955 -52387
rect 904 -22108 955 -22070
rect 904 -25161 955 -25123
rect 904 -47739 955 -47701
rect 904 -49159 955 -49121
rect 904 -64211 955 -64173
rect 904 -72376 955 -72338
rect 904 -36805 955 -36767
rect 904 -56259 955 -56221
rect 904 -15860 955 -15822
rect 904 -16783 955 -16745
rect 904 -23386 955 -23348
rect 904 -28924 955 -28886
rect 904 -13872 955 -13834
rect 904 -17138 955 -17100
rect 904 -9896 955 -9858
rect 904 -24664 955 -24626
rect 904 -12310 955 -12272
rect 904 -34817 955 -34779
rect 904 -66057 955 -66019
rect 904 -27220 955 -27182
rect 904 -16499 955 -16461
rect 904 -46745 955 -46707
rect 904 -66838 955 -66800
rect 904 -31267 955 -31229
rect 904 -34036 955 -33998
rect 904 -28285 955 -28247
rect 904 -19836 955 -19798
rect 904 -17706 955 -17668
rect 904 -12949 955 -12911
rect 904 -37657 955 -37619
rect 904 -34107 955 -34069
rect 904 -13020 955 -12982
rect 904 -53277 955 -53239
rect 904 -9115 955 -9077
rect 904 -16854 955 -16816
rect 904 -55407 955 -55369
rect 904 -51431 955 -51393
rect 904 -9186 955 -9148
rect 904 -64992 955 -64954
rect 904 -53135 955 -53097
rect 904 -26084 955 -26046
rect 904 -33255 955 -33217
rect 904 -71027 955 -70989
rect 904 -21540 955 -21502
rect 904 -18345 955 -18307
rect 904 -69678 955 -69640
rect 904 -33113 955 -33075
rect 904 -70175 955 -70137
rect 904 -30202 955 -30164
rect 904 -69607 955 -69569
rect 904 -11600 955 -11562
rect 904 -38367 955 -38329
rect 904 -55194 955 -55156
rect 904 -18913 955 -18875
rect 904 -20049 955 -20011
rect 904 -38793 955 -38755
rect 904 -64140 955 -64102
rect 904 -14653 955 -14615
rect 904 -22250 955 -22212
rect 904 -10606 955 -10568
rect 904 -21327 955 -21289
rect 904 -20262 955 -20224
rect 904 -12381 955 -12343
rect 904 -18842 955 -18804
rect 904 -11174 955 -11136
rect 904 -17919 955 -17881
rect 904 -10961 955 -10923
rect 904 -14085 955 -14047
rect 904 -69820 955 -69782
rect 904 -15931 955 -15893
rect 904 -67264 955 -67226
rect 904 -23812 955 -23774
rect 904 -37373 955 -37335
rect 904 -21256 955 -21218
rect 904 -18274 955 -18236
rect 904 -30557 955 -30519
rect 904 -22392 955 -22354
rect 904 -32119 955 -32081
rect 904 -14156 955 -14118
rect 904 -39787 955 -39749
rect 904 -12665 955 -12627
rect 904 -36521 955 -36483
rect 904 -11813 955 -11775
rect 904 -34888 955 -34850
rect 904 -55975 955 -55937
rect 904 -48307 955 -48269
rect 904 -13091 955 -13053
rect 904 -72305 955 -72267
rect 904 -22960 955 -22922
rect 904 -68329 955 -68291
rect 904 -35456 955 -35418
rect 904 -42059 955 -42021
rect 904 -59454 955 -59416
rect 904 -35243 955 -35205
rect 904 -30273 955 -30235
rect 904 -43621 955 -43583
rect 904 -52709 955 -52671
rect 904 -31906 955 -31868
rect 904 -54129 955 -54091
rect 904 -43337 955 -43299
rect 904 -49443 955 -49405
rect 904 -58673 955 -58635
rect 904 -43763 955 -43725
rect 904 -23528 955 -23490
rect 904 -11458 955 -11420
rect 904 -27149 955 -27111
rect 904 -17351 955 -17313
rect 904 -71240 955 -71202
rect 904 -61300 955 -61262
rect 904 -47029 955 -46991
rect 904 -28569 955 -28531
rect 904 -66625 955 -66587
rect 904 -58105 955 -58067
rect 904 -28356 955 -28318
rect 904 -19978 955 -19940
rect 904 -69465 955 -69427
rect 904 -34462 955 -34424
rect 904 -26439 955 -26401
rect 904 -27433 955 -27395
rect 904 -23883 955 -23845
rect 904 -12097 955 -12059
rect 904 -20120 955 -20082
rect 904 -14795 955 -14757
rect 904 -49869 955 -49831
rect 904 -63075 955 -63037
rect 904 -28001 955 -27963
rect 904 -11316 955 -11278
rect 904 -34533 955 -34495
rect 904 -72447 955 -72409
rect 904 -27007 955 -26969
rect 904 -25658 955 -25620
rect 904 -18487 955 -18449
rect 904 -33326 955 -33288
rect 904 -51147 955 -51109
rect 904 -20830 955 -20792
rect 904 -15647 955 -15609
rect 904 -29918 955 -29880
rect 904 -48875 955 -48837
rect 904 -13659 955 -13621
rect 904 -9967 955 -9929
rect 904 -54413 955 -54375
rect 904 -47597 955 -47559
rect 904 -29492 955 -29454
rect 904 -32829 955 -32791
rect 904 -33752 955 -33714
rect 904 -10038 955 -10000
rect 904 -30415 955 -30377
rect 904 -13162 955 -13124
rect 904 -26865 955 -26827
rect 904 -16002 955 -15964
rect 904 -38083 955 -38045
rect 904 -9399 955 -9361
rect 904 -51573 955 -51535
rect 904 -16996 955 -16958
rect 904 -12523 955 -12485
rect 904 -31480 955 -31442
rect 904 -20191 955 -20153
rect 904 -38225 955 -38187
rect 904 -21611 955 -21573
rect 904 -28711 955 -28673
rect 904 -26794 955 -26756
rect 904 -44331 955 -44293
rect 904 -44047 955 -44009
rect 904 -66412 955 -66374
rect 904 -23954 955 -23916
rect 904 -20972 955 -20934
rect 904 -17635 955 -17597
rect 904 -34391 955 -34353
rect 904 -13801 955 -13763
rect 904 -60448 955 -60410
rect 904 -42343 955 -42305
rect 904 -36237 955 -36199
rect 904 -12168 955 -12130
rect 904 -14582 955 -14544
rect 904 -46319 955 -46281
rect 904 -51999 955 -51961
rect 904 -42485 955 -42447
rect 904 -19765 955 -19727
rect 904 -20617 955 -20579
rect 904 -35811 955 -35773
rect 904 -63572 955 -63534
rect 904 -46603 955 -46565
rect 904 -44757 955 -44719
rect 904 -42769 955 -42731
rect 904 -71737 955 -71699
rect 904 -52993 955 -52955
rect 904 -56756 955 -56718
rect 904 -19339 955 -19301
rect 738 -36095 789 -36057
rect 738 -42911 789 -42873
rect 738 -10535 789 -10497
rect 738 -66980 789 -66942
rect 738 -51360 789 -51322
rect 738 -42627 789 -42589
rect 738 -15363 789 -15325
rect 738 -26013 789 -25975
rect 738 -34675 789 -34637
rect 738 -54200 789 -54162
rect 738 -20901 789 -20863
rect 738 -11245 789 -11207
rect 738 -28143 789 -28105
rect 738 -39432 789 -39394
rect 738 -31977 789 -31939
rect 738 -41420 789 -41382
rect 738 -43124 789 -43086
rect 738 -68116 789 -68078
rect 738 -48520 789 -48482
rect 738 -15008 789 -14970
rect 738 -68684 789 -68646
rect 738 -16144 789 -16106
rect 738 -10819 789 -10781
rect 738 -65347 789 -65309
rect 738 -43195 789 -43157
rect 738 -22463 789 -22425
rect 738 -9257 789 -9219
rect 738 -62933 789 -62895
rect 738 -13304 789 -13266
rect 738 -24451 789 -24413
rect 738 -43692 789 -43654
rect 738 -49727 789 -49689
rect 738 -10180 789 -10142
rect 738 -23457 789 -23419
rect 738 -11742 789 -11704
rect 738 -35527 789 -35489
rect 738 -16357 789 -16319
rect 738 -24025 789 -23987
rect 738 -25729 789 -25691
rect 738 -58602 789 -58564
rect 738 -20759 789 -20721
rect 738 -35953 789 -35915
rect 738 -66341 789 -66303
rect 738 -13517 789 -13479
rect 738 -49656 789 -49618
rect 738 -62365 789 -62327
rect 738 -17280 789 -17242
rect 738 -51076 789 -51038
rect 738 -43479 789 -43441
rect 738 -31551 789 -31513
rect 738 -22037 789 -21999
rect 738 -27291 789 -27253
rect 738 -58886 789 -58848
rect 738 -65986 789 -65948
rect 738 -72163 789 -72125
rect 738 -38935 789 -38897
rect 738 -52780 789 -52742
rect 738 -20333 789 -20295
rect 738 -15718 789 -15680
rect 738 -62862 789 -62824
rect 738 -52567 789 -52529
rect 738 -19055 789 -19017
rect 738 -43408 789 -43370
rect 738 -54271 789 -54233
rect 738 -61939 789 -61901
rect 738 -50579 789 -50541
rect 738 -67406 789 -67368
rect 738 -31693 789 -31655
rect 738 -42272 789 -42234
rect 738 -12594 789 -12556
rect 738 -26297 789 -26259
rect 738 -64353 789 -64315
rect 738 -14440 789 -14402
rect 738 -46035 789 -45997
rect 738 -66483 789 -66445
rect 738 -24877 789 -24839
rect 738 -28853 789 -28815
rect 738 -35385 789 -35347
rect 738 -40852 789 -40814
rect 738 -9683 789 -9645
rect 738 -56330 789 -56292
rect 738 -70956 789 -70918
rect 738 -10464 789 -10426
rect 738 -50863 789 -50825
rect 738 -59738 789 -59700
rect 738 -59170 789 -59132
rect 738 -15292 789 -15254
rect 738 -38651 789 -38613
rect 738 -12736 789 -12698
rect 738 -60803 789 -60765
rect 738 -30841 789 -30803
rect 738 -34959 789 -34921
rect 738 -42556 789 -42518
rect 738 -33397 789 -33359
rect 738 -47455 789 -47417
rect 738 -52283 789 -52245
rect 738 -29563 789 -29525
rect 738 -44615 789 -44577
rect 738 -32971 789 -32933
rect 738 -40355 789 -40317
rect 738 -45112 789 -45074
rect 738 -15576 789 -15538
rect 738 -60590 789 -60552
rect 738 -68755 789 -68717
rect 738 -46248 789 -46210
rect 738 -32687 789 -32649
rect 738 -66696 789 -66658
rect 738 -21753 789 -21715
rect 738 -17564 789 -17526
rect 738 -55762 789 -55724
rect 738 -65276 789 -65238
rect 738 -11032 789 -10994
rect 738 -58531 789 -58493
rect 738 -53064 789 -53026
rect 738 -14511 789 -14473
rect 738 -22605 789 -22567
rect 738 -55123 789 -55085
rect 738 -68471 789 -68433
rect 738 -65631 789 -65593
rect 738 -17990 789 -17952
rect 738 -29989 789 -29951
rect 738 -60377 789 -60339
rect 738 -63856 789 -63818
rect 738 -40284 789 -40246
rect 738 -11103 789 -11065
rect 738 -63288 789 -63250
rect 738 -14866 789 -14828
rect 738 -21469 789 -21431
rect 738 -23599 789 -23561
rect 738 -11884 789 -11846
rect 738 -55549 789 -55511
rect 738 -11529 789 -11491
rect 738 -15434 789 -15396
rect 738 -64069 789 -64031
rect 738 -32403 789 -32365
rect 738 -17209 789 -17171
rect 738 -51715 789 -51677
rect 738 -18771 789 -18733
rect 738 -25587 789 -25549
rect 738 -56117 789 -56079
rect 738 -51644 789 -51606
rect 738 -72092 789 -72054
rect 738 -9825 789 -9787
rect 738 -12807 789 -12769
rect 738 -21185 789 -21147
rect 738 -32261 789 -32223
rect 738 -33539 789 -33501
rect 738 -25019 789 -24981
rect 738 -63643 789 -63605
rect 738 -53916 789 -53878
rect 738 -19907 789 -19869
rect 738 -57466 789 -57428
rect 738 -18629 789 -18591
rect 738 -33681 789 -33643
rect 738 -10677 789 -10639
rect 738 -13588 789 -13550
rect 738 -22747 789 -22709
rect 738 -29847 789 -29809
rect 738 -48023 789 -47985
rect 738 -27717 789 -27679
rect 738 -62010 789 -61972
rect 738 -44899 789 -44861
rect 738 -49088 789 -49050
rect 738 -17422 789 -17384
rect 738 -47952 789 -47914
rect 738 -30131 789 -30093
rect 738 -45183 789 -45145
rect 738 -45467 789 -45429
rect 738 -23741 789 -23703
rect 738 -60306 789 -60268
rect 738 -24593 789 -24555
rect 738 -23173 789 -23135
rect 738 -14937 789 -14899
rect 738 -32545 789 -32507
rect 738 -20475 789 -20437
rect 738 -10890 789 -10852
rect 738 -18132 789 -18094
rect 738 -14724 789 -14686
rect 738 -10748 789 -10710
rect 738 -52212 789 -52174
rect 738 -12239 789 -12201
rect 738 -33965 789 -33927
rect 738 -37231 789 -37193
rect 738 -41775 789 -41737
rect 738 -50508 789 -50470
rect 738 -33823 789 -33785
rect 738 -41491 789 -41453
rect 738 -22179 789 -22141
rect 738 -24735 789 -24697
rect 738 -39503 789 -39465
rect 738 -19481 789 -19443
rect 738 -40071 789 -40033
rect 738 -21043 789 -21005
rect 738 -61371 789 -61333
rect 738 -10393 789 -10355
rect 738 -29705 789 -29667
rect 738 -31835 789 -31797
rect 738 -29279 789 -29241
rect 738 -9470 789 -9432
rect 738 -11671 789 -11633
rect 738 -60093 789 -60055
rect 738 -19197 789 -19159
rect 738 -13943 789 -13905
rect 738 -53419 789 -53381
rect 738 -64495 789 -64457
rect 738 -14298 789 -14260
rect 738 -65773 789 -65735
rect 738 -23315 789 -23277
rect 738 -35669 789 -35631
rect 738 -44544 789 -44506
rect 738 -25871 789 -25833
rect 738 -24167 789 -24129
rect 738 -29137 789 -29099
rect 738 -45751 789 -45713
rect 738 -59880 789 -59842
rect 738 -11955 789 -11917
rect 738 -37515 789 -37477
rect 738 -61016 789 -60978
rect 738 -63217 789 -63179
rect 738 -14014 789 -13976
rect 738 -17848 789 -17810
rect 738 -41136 789 -41098
rect 738 -68045 789 -68007
rect 738 -60022 789 -59984
rect 738 -69039 789 -69001
rect 738 -63927 789 -63889
rect 738 -14369 789 -14331
rect 738 -34249 789 -34211
rect 738 -24309 789 -24271
rect 738 -47171 789 -47133
rect 738 -28427 789 -28389
rect 738 -15150 789 -15112
rect 738 -15221 789 -15183
rect 738 -70530 789 -70492
rect 738 -69749 789 -69711
rect 738 -52496 789 -52458
rect 738 -47100 789 -47062
rect 738 -44260 789 -44222
rect 738 -69252 789 -69214
rect 738 -36947 789 -36909
rect 738 -16712 789 -16674
rect 738 -42840 789 -42802
rect 738 -50295 789 -50257
rect 738 -9328 789 -9290
rect 738 -12026 789 -11988
rect 738 -38012 789 -37974
rect 738 -9541 789 -9503
rect 738 -11387 789 -11349
rect 738 -71311 789 -71273
rect 738 -14227 789 -14189
rect 738 -26581 789 -26543
rect 738 -15505 789 -15467
rect 738 -16286 789 -16248
rect 738 -22889 789 -22851
rect 738 -63501 789 -63463
rect 738 -26723 789 -26685
rect 738 -16925 789 -16887
rect 738 -48591 789 -48553
rect 738 -37799 789 -37761
rect 738 -41207 789 -41169
rect 738 -40639 789 -40601
rect 738 -10251 789 -10213
rect 738 -60945 789 -60907
rect 738 -67548 789 -67510
rect 738 -64708 789 -64670
rect 738 -12878 789 -12840
rect 738 -36663 789 -36625
rect 738 -70672 789 -70634
rect 738 -63714 789 -63676
rect 738 -18061 789 -18023
rect 738 -9754 789 -9716
rect 738 -30699 789 -30661
rect 738 -55904 789 -55866
rect 738 -61158 789 -61120
rect 738 -53703 789 -53665
rect 738 -40923 789 -40885
rect 738 -36592 789 -36554
rect 738 -70317 789 -70279
rect 738 -56614 789 -56576
rect 738 -58247 789 -58209
rect 738 -16428 789 -16390
rect 738 -35101 789 -35063
rect 738 -50011 789 -49973
rect 738 -10109 789 -10071
rect 738 -13233 789 -13195
rect 738 -12452 789 -12414
rect 738 -13446 789 -13408
rect 738 -50224 789 -50186
rect 738 -57679 789 -57641
rect 738 -13375 789 -13337
rect 738 -65915 789 -65877
rect 738 -16641 789 -16603
rect 738 -50792 789 -50754
rect 738 -55691 789 -55653
rect 738 -16570 789 -16532
rect 738 -31409 789 -31371
rect 738 -17493 789 -17455
rect 738 -40000 789 -39962
rect 738 -45396 789 -45358
rect 738 -38864 789 -38826
rect 738 -27575 789 -27537
rect 738 -29421 789 -29383
rect 738 -46887 789 -46849
rect 738 -48236 789 -48198
rect 738 -53987 789 -53949
rect 738 -57963 789 -57925
rect 738 -44828 789 -44790
rect 738 -22321 789 -22283
rect 738 -15789 789 -15751
rect 738 -17067 789 -17029
rect 738 -40568 789 -40530
rect 738 -28995 789 -28957
rect 738 -52851 789 -52813
rect 738 -69323 789 -69285
rect 738 -47668 789 -47630
rect 738 -71169 789 -71131
rect 738 -26155 789 -26117
rect 738 -31125 789 -31087
rect 738 -37444 789 -37406
rect 738 -27859 789 -27821
rect 738 -15079 789 -15041
rect 738 -70814 789 -70776
rect 738 -25303 789 -25265
rect 738 -13730 789 -13692
rect 738 -23031 789 -22993
rect 738 -16215 789 -16177
rect 738 -25445 789 -25407
rect 738 -39219 789 -39181
rect 738 -19623 789 -19585
rect 738 -66128 789 -66090
rect 738 -56472 789 -56434
rect 738 -63430 789 -63392
rect 738 -16073 789 -16035
rect 738 -10322 789 -10284
rect 738 -41988 789 -41950
rect 738 -71595 789 -71557
rect 738 -55052 789 -55014
rect 738 -64921 789 -64883
rect 738 -45680 789 -45642
rect 738 -58815 789 -58777
rect 738 -71524 789 -71486
rect 738 -43976 789 -43938
rect 738 -65134 789 -65096
rect 738 -48804 789 -48766
rect 738 -57111 789 -57073
rect 738 -38296 789 -38258
rect 738 -49372 789 -49334
rect 738 -45964 789 -45926
rect 738 -21895 789 -21857
rect 738 -57750 789 -57712
rect 738 -9612 789 -9574
rect 738 -46532 789 -46494
rect 738 -67832 789 -67794
rect 738 -61797 789 -61759
rect 738 -63785 789 -63747
rect 738 -30983 789 -30945
rect 738 -17777 789 -17739
rect 738 -53348 789 -53310
rect 738 -49940 789 -49902
rect 738 -25161 789 -25123
rect 738 -47739 789 -47701
rect 738 -49159 789 -49121
rect 738 -62791 789 -62753
rect 738 -15860 789 -15822
rect 738 -16783 789 -16745
rect 738 -13872 789 -13834
rect 738 -17138 789 -17100
rect 738 -9896 789 -9858
rect 738 -12310 789 -12272
rect 738 -34817 789 -34779
rect 738 -16499 789 -16461
rect 738 -31267 789 -31229
rect 738 -28285 789 -28247
rect 738 -17706 789 -17668
rect 738 -12949 789 -12911
rect 738 -66909 789 -66871
rect 738 -34107 789 -34069
rect 738 -13020 789 -12982
rect 738 -9115 789 -9077
rect 738 -16854 789 -16816
rect 738 -51431 789 -51393
rect 738 -9186 789 -9148
rect 738 -53135 789 -53097
rect 738 -33255 789 -33217
rect 738 -18345 789 -18307
rect 738 -33113 789 -33075
rect 738 -70175 789 -70137
rect 738 -62578 789 -62540
rect 738 -69607 789 -69569
rect 738 -11600 789 -11562
rect 738 -38367 789 -38329
rect 738 -55194 789 -55156
rect 738 -18913 789 -18875
rect 738 -67761 789 -67723
rect 738 -20049 789 -20011
rect 738 -14653 789 -14615
rect 738 -63998 789 -63960
rect 738 -10606 789 -10568
rect 738 -21327 789 -21289
rect 738 -12381 789 -12343
rect 738 -11174 789 -11136
rect 738 -17919 789 -17881
rect 738 -10961 789 -10923
rect 738 -14085 789 -14047
rect 738 -63359 789 -63321
rect 738 -39148 789 -39110
rect 738 -69820 789 -69782
rect 738 -59241 789 -59203
rect 738 -15931 789 -15893
rect 738 -66270 789 -66232
rect 738 -67264 789 -67226
rect 738 -41704 789 -41666
rect 738 -62152 789 -62114
rect 738 -30557 789 -30519
rect 738 -36876 789 -36838
rect 738 -32119 789 -32081
rect 738 -14156 789 -14118
rect 738 -39787 789 -39749
rect 738 -12665 789 -12627
rect 738 -11813 789 -11775
rect 738 -55975 789 -55937
rect 738 -48307 789 -48269
rect 738 -67477 789 -67439
rect 738 -13091 789 -13053
rect 738 -68400 789 -68362
rect 738 -71808 789 -71770
rect 738 -42059 789 -42021
rect 738 -55478 789 -55440
rect 738 -59454 789 -59416
rect 738 -35243 789 -35205
rect 738 -30273 789 -30235
rect 738 -49443 789 -49405
rect 738 -43763 789 -43725
rect 738 -11458 789 -11420
rect 738 -27149 789 -27111
rect 738 -17351 789 -17313
rect 738 -61300 789 -61262
rect 738 -37160 789 -37122
rect 738 -69536 789 -69498
rect 738 -28569 789 -28531
rect 738 -69962 789 -69924
rect 738 -26439 789 -26401
rect 738 -56969 789 -56931
rect 738 -27433 789 -27395
rect 738 -23883 789 -23845
rect 738 -12097 789 -12059
rect 738 -14795 789 -14757
rect 738 -28001 789 -27963
rect 738 -11316 789 -11278
rect 738 -34533 789 -34495
rect 738 -61655 789 -61617
rect 738 -27007 789 -26969
rect 738 -61513 789 -61475
rect 738 -18487 789 -18449
rect 738 -59525 789 -59487
rect 738 -51147 789 -51109
rect 738 -46816 789 -46778
rect 738 -15647 789 -15609
rect 738 -48875 789 -48837
rect 738 -13659 789 -13621
rect 738 -9967 789 -9929
rect 738 -57537 789 -57499
rect 738 -57324 789 -57286
rect 738 -58034 789 -57996
rect 738 -32829 789 -32791
rect 738 -10038 789 -10000
rect 738 -30415 789 -30377
rect 738 -13162 789 -13124
rect 738 -26865 789 -26827
rect 738 -64424 789 -64386
rect 738 -16002 789 -15964
rect 738 -47384 789 -47346
rect 738 -38083 789 -38045
rect 738 -9399 789 -9361
rect 738 -16996 789 -16958
rect 738 -72234 789 -72196
rect 738 -51928 789 -51890
rect 738 -12523 789 -12485
rect 738 -20191 789 -20153
rect 738 -21611 789 -21573
rect 738 -28711 789 -28673
rect 738 -38580 789 -38542
rect 738 -37728 789 -37690
rect 738 -44331 789 -44293
rect 738 -44047 789 -44009
rect 738 -17635 789 -17597
rect 738 -59809 789 -59771
rect 738 -65489 789 -65451
rect 738 -34391 789 -34353
rect 738 -13801 789 -13763
rect 738 -71382 789 -71344
rect 738 -42343 789 -42305
rect 738 -53632 789 -53594
rect 738 -36237 789 -36199
rect 738 -12168 789 -12130
rect 738 -14582 789 -14544
rect 738 -46319 789 -46281
rect 738 -51999 789 -51961
rect 738 -39716 789 -39678
rect 738 -67193 789 -67155
rect 738 -19765 789 -19727
rect 738 -20617 789 -20579
rect 738 -35811 789 -35773
rect 738 -54484 789 -54446
rect 738 -63572 789 -63534
rect 738 -46603 789 -46565
rect 738 -71737 789 -71699
rect 738 -56756 789 -56718
rect 738 -19339 789 -19301
rect 655 -36095 706 -36057
rect 655 -29634 706 -29596
rect 655 -10535 706 -10497
rect 655 -42627 706 -42589
rect 655 -15363 706 -15325
rect 655 -34675 706 -34637
rect 655 -43053 706 -43015
rect 655 -11245 706 -11207
rect 655 -41349 706 -41311
rect 655 -71950 706 -71912
rect 655 -28143 706 -28105
rect 655 -31338 706 -31300
rect 655 -55265 706 -55227
rect 655 -56827 706 -56789
rect 655 -37941 706 -37903
rect 655 -41420 706 -41382
rect 655 -43124 706 -43086
rect 655 -70743 706 -70705
rect 655 -15008 706 -14970
rect 655 -16144 706 -16106
rect 655 -10819 706 -10781
rect 655 -59951 706 -59913
rect 655 -43195 706 -43157
rect 655 -22463 706 -22425
rect 655 -9257 706 -9219
rect 655 -13304 706 -13266
rect 655 -20688 706 -20650
rect 655 -24451 706 -24413
rect 655 -43692 706 -43654
rect 655 -10180 706 -10142
rect 655 -29350 706 -29312
rect 655 -11742 706 -11704
rect 655 -35527 706 -35489
rect 655 -16357 706 -16319
rect 655 -64850 706 -64812
rect 655 -20759 706 -20721
rect 655 -62436 706 -62398
rect 655 -13517 706 -13479
rect 655 -53845 706 -53807
rect 655 -17280 706 -17242
rect 655 -51076 706 -51038
rect 655 -31551 706 -31513
rect 655 -27291 706 -27253
rect 655 -58886 706 -58848
rect 655 -65986 706 -65948
rect 655 -52780 706 -52742
rect 655 -55336 706 -55298
rect 655 -51005 706 -50967
rect 655 -15718 706 -15680
rect 655 -19055 706 -19017
rect 655 -50579 706 -50541
rect 655 -50934 706 -50896
rect 655 -12594 706 -12556
rect 655 -45822 706 -45784
rect 655 -62507 706 -62469
rect 655 -14440 706 -14402
rect 655 -37302 706 -37264
rect 655 -46035 706 -45997
rect 655 -66483 706 -66445
rect 655 -27930 706 -27892
rect 655 -40852 706 -40814
rect 655 -9683 706 -9645
rect 655 -56330 706 -56292
rect 655 -70956 706 -70918
rect 655 -10464 706 -10426
rect 655 -42414 706 -42376
rect 655 -15292 706 -15254
rect 655 -46461 706 -46423
rect 655 -38651 706 -38613
rect 655 -41278 706 -41240
rect 655 -59028 706 -58990
rect 655 -12736 706 -12698
rect 655 -25516 706 -25478
rect 655 -34746 706 -34708
rect 655 -36166 706 -36128
rect 655 -35314 706 -35276
rect 655 -60803 706 -60765
rect 655 -34959 706 -34921
rect 655 -64282 706 -64244
rect 655 -42556 706 -42518
rect 655 -55833 706 -55795
rect 655 -52283 706 -52245
rect 655 -29563 706 -29525
rect 655 -40142 706 -40104
rect 655 -48733 706 -48695
rect 655 -69394 706 -69356
rect 655 -32971 706 -32933
rect 655 -40355 706 -40317
rect 655 -27646 706 -27608
rect 655 -15576 706 -15538
rect 655 -60590 706 -60552
rect 655 -41917 706 -41879
rect 655 -68755 706 -68717
rect 655 -32758 706 -32720
rect 655 -39645 706 -39607
rect 655 -32687 706 -32649
rect 655 -66696 706 -66658
rect 655 -17564 706 -17526
rect 655 -11032 706 -10994
rect 655 -63146 706 -63108
rect 655 -58531 706 -58493
rect 655 -38438 706 -38400
rect 655 -14511 706 -14473
rect 655 -68968 706 -68930
rect 655 -17990 706 -17952
rect 655 -32474 706 -32436
rect 655 -60377 706 -60339
rect 655 -35598 706 -35560
rect 655 -40284 706 -40246
rect 655 -63856 706 -63818
rect 655 -11103 706 -11065
rect 655 -63288 706 -63250
rect 655 -35882 706 -35844
rect 655 -14866 706 -14828
rect 655 -23599 706 -23561
rect 655 -62081 706 -62043
rect 655 -11884 706 -11846
rect 655 -55549 706 -55511
rect 655 -11529 706 -11491
rect 655 -15434 706 -15396
rect 655 -64069 706 -64031
rect 655 -32403 706 -32365
rect 655 -17209 706 -17171
rect 655 -51715 706 -51677
rect 655 -33894 706 -33856
rect 655 -18771 706 -18733
rect 655 -49230 706 -49192
rect 655 -25587 706 -25549
rect 655 -68613 706 -68575
rect 655 -51644 706 -51606
rect 655 -9825 706 -9787
rect 655 -52141 706 -52103
rect 655 -52638 706 -52600
rect 655 -70459 706 -70421
rect 655 -12807 706 -12769
rect 655 -44189 706 -44151
rect 655 -57040 706 -57002
rect 655 -33539 706 -33501
rect 655 -25019 706 -24981
rect 655 -40781 706 -40743
rect 655 -36734 706 -36696
rect 655 -63643 706 -63605
rect 655 -25232 706 -25194
rect 655 -53916 706 -53878
rect 655 -39077 706 -39039
rect 655 -56543 706 -56505
rect 655 -19907 706 -19869
rect 655 -26936 706 -26898
rect 655 -10677 706 -10639
rect 655 -65205 706 -65167
rect 655 -13588 706 -13550
rect 655 -22747 706 -22709
rect 655 -32190 706 -32152
rect 655 -29847 706 -29809
rect 655 -50437 706 -50399
rect 655 -71879 706 -71841
rect 655 -44899 706 -44861
rect 655 -66767 706 -66729
rect 655 -17422 706 -17384
rect 655 -24096 706 -24058
rect 655 -30131 706 -30093
rect 655 -45467 706 -45429
rect 655 -60164 706 -60126
rect 655 -29066 706 -29028
rect 655 -14937 706 -14899
rect 655 -20475 706 -20437
rect 655 -53774 706 -53736
rect 655 -10890 706 -10852
rect 655 -18132 706 -18094
rect 655 -14724 706 -14686
rect 655 -49301 706 -49263
rect 655 -10748 706 -10710
rect 655 -33610 706 -33572
rect 655 -52212 706 -52174
rect 655 -12239 706 -12201
rect 655 -24380 706 -24342
rect 655 -50508 706 -50470
rect 655 -49798 706 -49760
rect 655 -19268 706 -19230
rect 655 -33823 706 -33785
rect 655 -41491 706 -41453
rect 655 -18416 706 -18378
rect 655 -60519 706 -60481
rect 655 -47526 706 -47488
rect 655 -68258 706 -68220
rect 655 -22179 706 -22141
rect 655 -24735 706 -24697
rect 655 -26652 706 -26614
rect 655 -23244 706 -23206
rect 655 -21043 706 -21005
rect 655 -10393 706 -10355
rect 655 -26368 706 -26330
rect 655 -31835 706 -31797
rect 655 -29279 706 -29241
rect 655 -9470 706 -9432
rect 655 -11671 706 -11633
rect 655 -46958 706 -46920
rect 655 -48165 706 -48127
rect 655 -13943 706 -13905
rect 655 -53419 706 -53381
rect 655 -30770 706 -30732
rect 655 -14298 706 -14260
rect 655 -65773 706 -65735
rect 655 -51502 706 -51464
rect 655 -23315 706 -23277
rect 655 -31622 706 -31584
rect 655 -25871 706 -25833
rect 655 -24167 706 -24129
rect 655 -11955 706 -11917
rect 655 -37515 706 -37477
rect 655 -59596 706 -59558
rect 655 -61016 706 -60978
rect 655 -63217 706 -63179
rect 655 -14014 706 -13976
rect 655 -22676 706 -22638
rect 655 -38509 706 -38471
rect 655 -17848 706 -17810
rect 655 -35030 706 -34992
rect 655 -60732 706 -60694
rect 655 -68045 706 -68007
rect 655 -60022 706 -59984
rect 655 -63927 706 -63889
rect 655 -14369 706 -14331
rect 655 -47171 706 -47133
rect 655 -28427 706 -28389
rect 655 -15150 706 -15112
rect 655 -15221 706 -15183
rect 655 -25800 706 -25762
rect 655 -69749 706 -69711
rect 655 -47100 706 -47062
rect 655 -44260 706 -44222
rect 655 -71453 706 -71415
rect 655 -36947 706 -36909
rect 655 -16712 706 -16674
rect 655 -58318 706 -58280
rect 655 -9328 706 -9290
rect 655 -12026 706 -11988
rect 655 -18984 706 -18946
rect 655 -38012 706 -37974
rect 655 -33042 706 -33004
rect 655 -9541 706 -9503
rect 655 -11387 706 -11349
rect 655 -71311 706 -71273
rect 655 -14227 706 -14189
rect 655 -15505 706 -15467
rect 655 -16286 706 -16248
rect 655 -63501 706 -63463
rect 655 -26723 706 -26685
rect 655 -16925 706 -16887
rect 655 -10251 706 -10213
rect 655 -40213 706 -40175
rect 655 -64708 706 -64670
rect 655 -34178 706 -34140
rect 655 -12878 706 -12840
rect 655 -70672 706 -70634
rect 655 -63714 706 -63676
rect 655 -18061 706 -18023
rect 655 -9754 706 -9716
rect 655 -21824 706 -21786
rect 655 -30699 706 -30661
rect 655 -45893 706 -45855
rect 655 -55904 706 -55866
rect 655 -40923 706 -40885
rect 655 -56614 706 -56576
rect 655 -16428 706 -16390
rect 655 -50011 706 -49973
rect 655 -10109 706 -10071
rect 655 -13233 706 -13195
rect 655 -12452 706 -12414
rect 655 -13446 706 -13408
rect 655 -13375 706 -13337
rect 655 -16641 706 -16603
rect 655 -16570 706 -16532
rect 655 -17493 706 -17455
rect 655 -64779 706 -64741
rect 655 -72021 706 -71983
rect 655 -45396 706 -45358
rect 655 -27575 706 -27537
rect 655 -52070 706 -52032
rect 655 -68826 706 -68788
rect 655 -56188 706 -56150
rect 655 -39006 706 -38968
rect 655 -48236 706 -48198
rect 655 -53987 706 -53949
rect 655 -57963 706 -57925
rect 655 -58460 706 -58422
rect 655 -44686 706 -44648
rect 655 -30486 706 -30448
rect 655 -45325 706 -45287
rect 655 -44828 706 -44790
rect 655 -15789 706 -15751
rect 655 -17067 706 -17029
rect 655 -71098 706 -71060
rect 655 -28995 706 -28957
rect 655 -52851 706 -52813
rect 655 -69323 706 -69285
rect 655 -20404 706 -20366
rect 655 -70246 706 -70208
rect 655 -47668 706 -47630
rect 655 -24948 706 -24910
rect 655 -26155 706 -26117
rect 655 -37444 706 -37406
rect 655 -28214 706 -28176
rect 655 -53206 706 -53168
rect 655 -27859 706 -27821
rect 655 -15079 706 -15041
rect 655 -25303 706 -25265
rect 655 -13730 706 -13692
rect 655 -23031 706 -22993
rect 655 -27362 706 -27324
rect 655 -61726 706 -61688
rect 655 -65844 706 -65806
rect 655 -16215 706 -16177
rect 655 -59383 706 -59345
rect 655 -41846 706 -41808
rect 655 -19552 706 -19514
rect 655 -28782 706 -28744
rect 655 -39219 706 -39181
rect 655 -19623 706 -19585
rect 655 -63430 706 -63392
rect 655 -16073 706 -16035
rect 655 -10322 706 -10284
rect 655 -41988 706 -41950
rect 655 -18700 706 -18662
rect 655 -28498 706 -28460
rect 655 -31054 706 -31016
rect 655 -65134 706 -65096
rect 655 -67335 706 -67297
rect 655 -48804 706 -48766
rect 655 -57111 706 -57073
rect 655 -61229 706 -61191
rect 655 -49372 706 -49334
rect 655 -67690 706 -67652
rect 655 -45964 706 -45926
rect 655 -21895 706 -21857
rect 655 -57750 706 -57712
rect 655 -9612 706 -9574
rect 655 -69181 706 -69143
rect 655 -46532 706 -46494
rect 655 -67122 706 -67084
rect 655 -61797 706 -61759
rect 655 -67832 706 -67794
rect 655 -63785 706 -63747
rect 655 -30983 706 -30945
rect 655 -17777 706 -17739
rect 655 -46390 706 -46352
rect 655 -22108 706 -22070
rect 655 -53348 706 -53310
rect 655 -49940 706 -49902
rect 655 -47739 706 -47701
rect 655 -64211 706 -64173
rect 655 -36805 706 -36767
rect 655 -56259 706 -56221
rect 655 -15860 706 -15822
rect 655 -16783 706 -16745
rect 655 -13872 706 -13834
rect 655 -17138 706 -17100
rect 655 -9896 706 -9858
rect 655 -24664 706 -24626
rect 655 -39574 706 -39536
rect 655 -12310 706 -12272
rect 655 -66057 706 -66019
rect 655 -27220 706 -27182
rect 655 -16499 706 -16461
rect 655 -70033 706 -69995
rect 655 -31267 706 -31229
rect 655 -19836 706 -19798
rect 655 -44118 706 -44080
rect 655 -17706 706 -17668
rect 655 -12949 706 -12911
rect 655 -66909 706 -66871
rect 655 -34107 706 -34069
rect 655 -13020 706 -12982
rect 655 -53277 706 -53239
rect 655 -9115 706 -9077
rect 655 -16854 706 -16816
rect 655 -55407 706 -55369
rect 655 -9186 706 -9148
rect 655 -26084 706 -26046
rect 655 -33255 706 -33217
rect 655 -71027 706 -70989
rect 655 -21540 706 -21502
rect 655 -70175 706 -70137
rect 655 -30202 706 -30164
rect 655 -62578 706 -62540
rect 655 -11600 706 -11562
rect 655 -64140 706 -64102
rect 655 -14653 706 -14615
rect 655 -63998 706 -63960
rect 655 -10606 706 -10568
rect 655 -21327 706 -21289
rect 655 -12381 706 -12343
rect 655 -11174 706 -11136
rect 655 -17919 706 -17881
rect 655 -10961 706 -10923
rect 655 -14085 706 -14047
rect 655 -63359 706 -63321
rect 655 -57892 706 -57854
rect 655 -39148 706 -39110
rect 655 -40710 706 -40672
rect 655 -42982 706 -42944
rect 655 -59241 706 -59203
rect 655 -15931 706 -15893
rect 655 -66270 706 -66232
rect 655 -67264 706 -67226
rect 655 -23812 706 -23774
rect 655 -37373 706 -37335
rect 655 -62152 706 -62114
rect 655 -21256 706 -21218
rect 655 -36876 706 -36838
rect 655 -22392 706 -22354
rect 655 -32119 706 -32081
rect 655 -45254 706 -45216
rect 655 -67903 706 -67865
rect 655 -48094 706 -48056
rect 655 -14156 706 -14118
rect 655 -39787 706 -39749
rect 655 -12665 706 -12627
rect 655 -11813 706 -11775
rect 655 -55975 706 -55937
rect 655 -48307 706 -48269
rect 655 -67477 706 -67439
rect 655 -13091 706 -13053
rect 655 -22960 706 -22922
rect 655 -68400 706 -68362
rect 655 -71808 706 -71770
rect 655 -48662 706 -48624
rect 655 -42059 706 -42021
rect 655 -55478 706 -55440
rect 655 -59454 706 -59416
rect 655 -35243 706 -35205
rect 655 -43621 706 -43583
rect 655 -52709 706 -52671
rect 655 -31906 706 -31868
rect 655 -49443 706 -49405
rect 655 -58673 706 -58635
rect 655 -43763 706 -43725
rect 655 -23528 706 -23490
rect 655 -11458 706 -11420
rect 655 -17351 706 -17313
rect 655 -61300 706 -61262
rect 655 -47029 706 -46991
rect 655 -43550 706 -43512
rect 655 -37870 706 -37832
rect 655 -69536 706 -69498
rect 655 -69962 706 -69924
rect 655 -58105 706 -58067
rect 655 -63004 706 -62966
rect 655 -34462 706 -34424
rect 655 -26439 706 -26401
rect 655 -50366 706 -50328
rect 655 -65560 706 -65522
rect 655 -54342 706 -54304
rect 655 -23883 706 -23845
rect 655 -12097 706 -12059
rect 655 -20120 706 -20082
rect 655 -14795 706 -14757
rect 655 -49869 706 -49831
rect 655 -63075 706 -63037
rect 655 -11316 706 -11278
rect 655 -27007 706 -26969
rect 655 -61513 706 -61475
rect 655 -18487 706 -18449
rect 655 -33326 706 -33288
rect 655 -51147 706 -51109
rect 655 -61442 706 -61404
rect 655 -15647 706 -15609
rect 655 -29918 706 -29880
rect 655 -48875 706 -48837
rect 655 -57253 706 -57215
rect 655 -13659 706 -13621
rect 655 -9967 706 -9929
rect 655 -54413 706 -54375
rect 655 -47597 706 -47559
rect 655 -57537 706 -57499
rect 655 -57324 706 -57286
rect 655 -10038 706 -10000
rect 655 -30415 706 -30377
rect 655 -13162 706 -13124
rect 655 -16002 706 -15964
rect 655 -38083 706 -38045
rect 655 -9399 706 -9361
rect 655 -51573 706 -51535
rect 655 -16996 706 -16958
rect 655 -12523 706 -12485
rect 655 -20191 706 -20153
rect 655 -21611 706 -21573
rect 655 -28711 706 -28673
rect 655 -38580 706 -38542
rect 655 -44331 706 -44293
rect 655 -66554 706 -66516
rect 655 -20972 706 -20934
rect 655 -17635 706 -17597
rect 655 -59809 706 -59771
rect 655 -65489 706 -65451
rect 655 -34391 706 -34353
rect 655 -13801 706 -13763
rect 655 -71382 706 -71344
rect 655 -12168 706 -12130
rect 655 -14582 706 -14544
rect 655 -39716 706 -39678
rect 655 -42485 706 -42447
rect 655 -35811 706 -35773
rect 655 -54484 706 -54446
rect 655 -63572 706 -63534
rect 655 -46603 706 -46565
rect 655 -44757 706 -44719
rect 655 -71737 706 -71699
rect 655 -19339 706 -19301
rect 489 -29208 540 -29170
rect 489 -29634 540 -29596
rect 489 -10535 540 -10497
rect 489 -42911 540 -42873
rect 489 -15363 540 -15325
rect 489 -26013 540 -25975
rect 489 -34675 540 -34637
rect 489 -41633 540 -41595
rect 489 -20901 540 -20863
rect 489 -54200 540 -54162
rect 489 -43053 540 -43015
rect 489 -11245 540 -11207
rect 489 -39432 540 -39394
rect 489 -31338 540 -31300
rect 489 -31977 540 -31939
rect 489 -43124 540 -43086
rect 489 -48520 540 -48482
rect 489 -15008 540 -14970
rect 489 -68684 540 -68646
rect 489 -70743 540 -70705
rect 489 -16144 540 -16106
rect 489 -10819 540 -10781
rect 489 -65347 540 -65309
rect 489 -43195 540 -43157
rect 489 -24806 540 -24768
rect 489 -9257 540 -9219
rect 489 -62933 540 -62895
rect 489 -58957 540 -58919
rect 489 -13304 540 -13266
rect 489 -33184 540 -33146
rect 489 -67974 540 -67936
rect 489 -24451 540 -24413
rect 489 -49727 540 -49689
rect 489 -10180 540 -10142
rect 489 -57395 540 -57357
rect 489 -25374 540 -25336
rect 489 -11742 540 -11704
rect 489 -16357 540 -16319
rect 489 -58602 540 -58564
rect 489 -35953 540 -35915
rect 489 -66341 540 -66303
rect 489 -13517 540 -13479
rect 489 -49656 540 -49618
rect 489 -58176 540 -58138
rect 489 -17280 540 -17242
rect 489 -70388 540 -70350
rect 489 -49585 540 -49547
rect 489 -51076 540 -51038
rect 489 -22037 540 -21999
rect 489 -27291 540 -27253
rect 489 -47313 540 -47275
rect 489 -28072 540 -28034
rect 489 -20333 540 -20295
rect 489 -51005 540 -50967
rect 489 -15718 540 -15680
rect 489 -62862 540 -62824
rect 489 -54271 540 -54233
rect 489 -61939 540 -61901
rect 489 -43905 540 -43867
rect 489 -70885 540 -70847
rect 489 -50934 540 -50896
rect 489 -12594 540 -12556
rect 489 -19694 540 -19656
rect 489 -64353 540 -64315
rect 489 -14440 540 -14402
rect 489 -37302 540 -37264
rect 489 -24877 540 -24839
rect 489 -27930 540 -27892
rect 489 -35385 540 -35347
rect 489 -40852 540 -40814
rect 489 -9683 540 -9645
rect 489 -10464 540 -10426
rect 489 -50863 540 -50825
rect 489 -59738 540 -59700
rect 489 -60874 540 -60836
rect 489 -15292 540 -15254
rect 489 -46461 540 -46423
rect 489 -38651 540 -38613
rect 489 -59028 540 -58990
rect 489 -12736 540 -12698
rect 489 -46177 540 -46139
rect 489 -25516 540 -25478
rect 489 -34746 540 -34708
rect 489 -35314 540 -35276
rect 489 -26510 540 -26472
rect 489 -30841 540 -30803
rect 489 -64282 540 -64244
rect 489 -55833 540 -55795
rect 489 -47455 540 -47417
rect 489 -52283 540 -52245
rect 489 -29563 540 -29525
rect 489 -48733 540 -48695
rect 489 -69394 540 -69356
rect 489 -32971 540 -32933
rect 489 -45112 540 -45074
rect 489 -15576 540 -15538
rect 489 -60590 540 -60552
rect 489 -41917 540 -41879
rect 489 -29776 540 -29738
rect 489 -46248 540 -46210
rect 489 -67619 540 -67581
rect 489 -39645 540 -39607
rect 489 -50721 540 -50683
rect 489 -66696 540 -66658
rect 489 -17564 540 -17526
rect 489 -55762 540 -55724
rect 489 -65276 540 -65238
rect 489 -11032 540 -10994
rect 489 -63146 540 -63108
rect 489 -53064 540 -53026
rect 489 -38438 540 -38400
rect 489 -30912 540 -30874
rect 489 -14511 540 -14473
rect 489 -22605 540 -22567
rect 489 -21966 540 -21928
rect 489 -68968 540 -68930
rect 489 -17990 540 -17952
rect 489 -27504 540 -27466
rect 489 -32474 540 -32436
rect 489 -62720 540 -62682
rect 489 -63856 540 -63818
rect 489 -11103 540 -11065
rect 489 -44970 540 -44932
rect 489 -63288 540 -63250
rect 489 -35882 540 -35844
rect 489 -14866 540 -14828
rect 489 -21469 540 -21431
rect 489 -62081 540 -62043
rect 489 -11884 540 -11846
rect 489 -55620 540 -55582
rect 489 -11529 540 -11491
rect 489 -15434 540 -15396
rect 489 -64069 540 -64031
rect 489 -32403 540 -32365
rect 489 -17209 540 -17171
rect 489 -42698 540 -42660
rect 489 -48449 540 -48411
rect 489 -62649 540 -62611
rect 489 -18771 540 -18733
rect 489 -25587 540 -25549
rect 489 -68613 540 -68575
rect 489 -9825 540 -9787
rect 489 -52141 540 -52103
rect 489 -19126 540 -19088
rect 489 -12807 540 -12769
rect 489 -44189 540 -44151
rect 489 -57040 540 -57002
rect 489 -33539 540 -33501
rect 489 -25019 540 -24981
rect 489 -40781 540 -40743
rect 489 -63643 540 -63605
rect 489 -64637 540 -64599
rect 489 -56543 540 -56505
rect 489 -19907 540 -19869
rect 489 -57466 540 -57428
rect 489 -18629 540 -18591
rect 489 -33681 540 -33643
rect 489 -10677 540 -10639
rect 489 -65205 540 -65167
rect 489 -13588 540 -13550
rect 489 -22747 540 -22709
rect 489 -62010 540 -61972
rect 489 -21398 540 -21360
rect 489 -66767 540 -66729
rect 489 -40497 540 -40459
rect 489 -17422 540 -17384
rect 489 -30131 540 -30093
rect 489 -22534 540 -22496
rect 489 -45183 540 -45145
rect 489 -45467 540 -45429
rect 489 -60164 540 -60126
rect 489 -28640 540 -28602
rect 489 -40426 540 -40388
rect 489 -23741 540 -23703
rect 489 -29066 540 -29028
rect 489 -23173 540 -23135
rect 489 -14937 540 -14899
rect 489 -32545 540 -32507
rect 489 -20475 540 -20437
rect 489 -10890 540 -10852
rect 489 -18132 540 -18094
rect 489 -14724 540 -14686
rect 489 -10748 540 -10710
rect 489 -33610 540 -33572
rect 489 -52212 540 -52174
rect 489 -12239 540 -12201
rect 489 -24380 540 -24342
rect 489 -37231 540 -37193
rect 489 -41775 540 -41737
rect 489 -49798 540 -49760
rect 489 -19268 540 -19230
rect 489 -60519 540 -60481
rect 489 -47526 540 -47488
rect 489 -68258 540 -68220
rect 489 -22179 540 -22141
rect 489 -69891 540 -69853
rect 489 -39503 540 -39465
rect 489 -26652 540 -26614
rect 489 -23244 540 -23206
rect 489 -21043 540 -21005
rect 489 -61371 540 -61333
rect 489 -10393 540 -10355
rect 489 -29705 540 -29667
rect 489 -31835 540 -31797
rect 489 -9470 540 -9432
rect 489 -11671 540 -11633
rect 489 -60093 540 -60055
rect 489 -19197 540 -19159
rect 489 -13943 540 -13905
rect 489 -53419 540 -53381
rect 489 -64495 540 -64457
rect 489 -30770 540 -30732
rect 489 -14298 540 -14260
rect 489 -65773 540 -65735
rect 489 -23315 540 -23277
rect 489 -32048 540 -32010
rect 489 -27078 540 -27040
rect 489 -29137 540 -29099
rect 489 -39290 540 -39252
rect 489 -11955 540 -11917
rect 489 -37515 540 -37477
rect 489 -61016 540 -60978
rect 489 -50650 540 -50612
rect 489 -63217 540 -63179
rect 489 -14014 540 -13976
rect 489 -22676 540 -22638
rect 489 -38509 540 -38471
rect 489 -17848 540 -17810
rect 489 -56898 540 -56860
rect 489 -69039 540 -69001
rect 489 -63927 540 -63889
rect 489 -14369 540 -14331
rect 489 -34249 540 -34211
rect 489 -24309 540 -24271
rect 489 -28427 540 -28389
rect 489 -15150 540 -15112
rect 489 -15221 540 -15183
rect 489 -59312 540 -59274
rect 489 -69749 540 -69711
rect 489 -56401 540 -56363
rect 489 -44260 540 -44222
rect 489 -71453 540 -71415
rect 489 -16712 540 -16674
rect 489 -58318 540 -58280
rect 489 -42840 540 -42802
rect 489 -9328 540 -9290
rect 489 -12026 540 -11988
rect 489 -52922 540 -52884
rect 489 -33042 540 -33004
rect 489 -9541 540 -9503
rect 489 -11387 540 -11349
rect 489 -71311 540 -71273
rect 489 -64566 540 -64528
rect 489 -14227 540 -14189
rect 489 -24238 540 -24200
rect 489 -26581 540 -26543
rect 489 -15505 540 -15467
rect 489 -45041 540 -45003
rect 489 -18558 540 -18520
rect 489 -65418 540 -65380
rect 489 -16286 540 -16248
rect 489 -63501 540 -63463
rect 489 -26723 540 -26685
rect 489 -16925 540 -16887
rect 489 -48591 540 -48553
rect 489 -71666 540 -71628
rect 489 -40639 540 -40601
rect 489 -10251 540 -10213
rect 489 -60945 540 -60907
rect 489 -67548 540 -67510
rect 489 -34178 540 -34140
rect 489 -12878 540 -12840
rect 489 -70672 540 -70634
rect 489 -63714 540 -63676
rect 489 -18061 540 -18023
rect 489 -9754 540 -9716
rect 489 -30699 540 -30661
rect 489 -55904 540 -55866
rect 489 -25942 540 -25904
rect 489 -40923 540 -40885
rect 489 -70317 540 -70279
rect 489 -56614 540 -56576
rect 489 -58247 540 -58209
rect 489 -16428 540 -16390
rect 489 -50011 540 -49973
rect 489 -10109 540 -10071
rect 489 -13233 540 -13195
rect 489 -12452 540 -12414
rect 489 -13446 540 -13408
rect 489 -13375 540 -13337
rect 489 -34320 540 -34282
rect 489 -16641 540 -16603
rect 489 -65915 540 -65877
rect 489 -50792 540 -50754
rect 489 -55691 540 -55653
rect 489 -16570 540 -16532
rect 489 -31409 540 -31371
rect 489 -37018 540 -36980
rect 489 -17493 540 -17455
rect 489 -48378 540 -48340
rect 489 -23102 540 -23064
rect 489 -45396 540 -45358
rect 489 -52070 540 -52032
rect 489 -57963 540 -57925
rect 489 -36024 540 -35986
rect 489 -49514 540 -49476
rect 489 -45325 540 -45287
rect 489 -15789 540 -15751
rect 489 -17067 540 -17029
rect 489 -40568 540 -40530
rect 489 -28995 540 -28957
rect 489 -23670 540 -23632
rect 489 -30344 540 -30306
rect 489 -69323 540 -69285
rect 489 -20404 540 -20366
rect 489 -70246 540 -70208
rect 489 -47668 540 -47630
rect 489 -24948 540 -24910
rect 489 -26155 540 -26117
rect 489 -37444 540 -37406
rect 489 -53206 540 -53168
rect 489 -32616 540 -32578
rect 489 -27859 540 -27821
rect 489 -15079 540 -15041
rect 489 -70814 540 -70776
rect 489 -13730 540 -13692
rect 489 -54058 540 -54020
rect 489 -61868 540 -61830
rect 489 -27362 540 -27324
rect 489 -65844 540 -65806
rect 489 -39361 540 -39323
rect 489 -16215 540 -16177
rect 489 -59383 540 -59345
rect 489 -41846 540 -41808
rect 489 -25445 540 -25407
rect 489 -37089 540 -37051
rect 489 -57821 540 -57783
rect 489 -38154 540 -38116
rect 489 -51857 540 -51819
rect 489 -56472 540 -56434
rect 489 -63430 540 -63392
rect 489 -16073 540 -16035
rect 489 -10322 540 -10284
rect 489 -41988 540 -41950
rect 489 -71595 540 -71557
rect 489 -18700 540 -18662
rect 489 -28498 540 -28460
rect 489 -71524 540 -71486
rect 489 -43976 540 -43938
rect 489 -65134 540 -65096
rect 489 -48804 540 -48766
rect 489 -57111 540 -57073
rect 489 -38296 540 -38258
rect 489 -9612 540 -9574
rect 489 -46532 540 -46494
rect 489 -67122 540 -67084
rect 489 -67832 540 -67794
rect 489 -63785 540 -63747
rect 489 -17777 540 -17739
rect 489 -46390 540 -46352
rect 489 -22108 540 -22070
rect 489 -53348 540 -53310
rect 489 -49940 540 -49902
rect 489 -47739 540 -47701
rect 489 -64211 540 -64173
rect 489 -62791 540 -62753
rect 489 -15860 540 -15822
rect 489 -16783 540 -16745
rect 489 -13872 540 -13834
rect 489 -17138 540 -17100
rect 489 -9896 540 -9858
rect 489 -39574 540 -39536
rect 489 -12310 540 -12272
rect 489 -34817 540 -34779
rect 489 -27220 540 -27182
rect 489 -16499 540 -16461
rect 489 -66838 540 -66800
rect 489 -31267 540 -31229
rect 489 -47242 540 -47204
rect 489 -19836 540 -19798
rect 489 -44118 540 -44080
rect 489 -17706 540 -17668
rect 489 -12949 540 -12911
rect 489 -41562 540 -41524
rect 489 -34107 540 -34069
rect 489 -13020 540 -12982
rect 489 -53277 540 -53239
rect 489 -9115 540 -9077
rect 489 -46106 540 -46068
rect 489 -16854 540 -16816
rect 489 -9186 540 -9148
rect 489 -53135 540 -53097
rect 489 -26084 540 -26046
rect 489 -21540 540 -21502
rect 489 -33113 540 -33075
rect 489 -70175 540 -70137
rect 489 -30202 540 -30164
rect 489 -11600 540 -11562
rect 489 -38367 540 -38329
rect 489 -64140 540 -64102
rect 489 -14653 540 -14615
rect 489 -63998 540 -63960
rect 489 -10606 540 -10568
rect 489 -20262 540 -20224
rect 489 -12381 540 -12343
rect 489 -11174 540 -11136
rect 489 -17919 540 -17881
rect 489 -10961 540 -10923
rect 489 -14085 540 -14047
rect 489 -63359 540 -63321
rect 489 -57892 540 -57854
rect 489 -69110 540 -69072
rect 489 -69820 540 -69782
rect 489 -40710 540 -40672
rect 489 -42982 540 -42944
rect 489 -15931 540 -15893
rect 489 -66270 540 -66232
rect 489 -23812 540 -23774
rect 489 -37373 540 -37335
rect 489 -41704 540 -41666
rect 489 -62152 540 -62114
rect 489 -45254 540 -45216
rect 489 -67903 540 -67865
rect 489 -14156 540 -14118
rect 489 -39787 540 -39749
rect 489 -12665 540 -12627
rect 489 -11813 540 -11775
rect 489 -34888 540 -34850
rect 489 -55975 540 -55937
rect 489 -67477 540 -67439
rect 489 -13091 540 -13053
rect 489 -68329 540 -68291
rect 489 -35456 540 -35418
rect 489 -48662 540 -48624
rect 489 -42059 540 -42021
rect 489 -59454 540 -59416
rect 489 -35243 540 -35205
rect 489 -30273 540 -30235
rect 489 -31906 540 -31868
rect 489 -54129 540 -54091
rect 489 -58673 540 -58635
rect 489 -11458 540 -11420
rect 489 -27149 540 -27111
rect 489 -17351 540 -17313
rect 489 -37160 540 -37122
rect 489 -28569 540 -28531
rect 489 -63004 540 -62966
rect 489 -69465 540 -69427
rect 489 -56969 540 -56931
rect 489 -27433 540 -27395
rect 489 -54342 540 -54304
rect 489 -23883 540 -23845
rect 489 -12097 540 -12059
rect 489 -14795 540 -14757
rect 489 -49869 540 -49831
rect 489 -63075 540 -63037
rect 489 -28001 540 -27963
rect 489 -11316 540 -11278
rect 489 -61513 540 -61475
rect 489 -51147 540 -51109
rect 489 -20830 540 -20792
rect 489 -61442 540 -61404
rect 489 -15647 540 -15609
rect 489 -59667 540 -59629
rect 489 -48875 540 -48837
rect 489 -43834 540 -43796
rect 489 -13659 540 -13621
rect 489 -9967 540 -9929
rect 489 -54413 540 -54375
rect 489 -47597 540 -47559
rect 489 -57537 540 -57499
rect 489 -33752 540 -33714
rect 489 -10038 540 -10000
rect 489 -13162 540 -13124
rect 489 -64424 540 -64386
rect 489 -16002 540 -15964
rect 489 -47384 540 -47346
rect 489 -9399 540 -9361
rect 489 -16996 540 -16958
rect 489 -51928 540 -51890
rect 489 -12523 540 -12485
rect 489 -31480 540 -31442
rect 489 -38225 540 -38187
rect 489 -21611 540 -21573
rect 489 -38580 540 -38542
rect 489 -44331 540 -44293
rect 489 -44047 540 -44009
rect 489 -66412 540 -66374
rect 489 -20972 540 -20934
rect 489 -17635 540 -17597
rect 489 -59809 540 -59771
rect 489 -13801 540 -13763
rect 489 -71382 540 -71344
rect 489 -60448 540 -60410
rect 489 -12168 540 -12130
rect 489 -14582 540 -14544
rect 489 -46319 540 -46281
rect 489 -51999 540 -51961
rect 489 -39716 540 -39678
rect 489 -67193 540 -67155
rect 489 -19765 540 -19727
rect 489 -35811 540 -35773
rect 489 -54484 540 -54446
rect 489 -51786 540 -51748
rect 489 -63572 540 -63534
rect 489 -46603 540 -46565
rect 489 -42769 540 -42731
rect 489 -52993 540 -52955
rect 489 -19339 540 -19301
rect 406 -29634 457 -29596
rect 406 -42911 457 -42873
rect 406 -10535 457 -10497
rect 406 -66980 457 -66942
rect 406 -51360 457 -51322
rect 406 -42627 457 -42589
rect 406 -15363 457 -15325
rect 406 -26013 457 -25975
rect 406 -53490 457 -53452
rect 406 -54200 457 -54162
rect 406 -57182 457 -57144
rect 406 -43053 457 -43015
rect 406 -11245 457 -11207
rect 406 -37941 457 -37903
rect 406 -31977 457 -31939
rect 406 -43124 457 -43086
rect 406 -27788 457 -27750
rect 406 -15008 457 -14970
rect 406 -70743 457 -70705
rect 406 -16144 457 -16106
rect 406 -10819 457 -10781
rect 406 -43195 457 -43157
rect 406 -24806 457 -24768
rect 406 -51218 457 -51180
rect 406 -22463 457 -22425
rect 406 -9257 457 -9219
rect 406 -62933 457 -62895
rect 406 -58957 457 -58919
rect 406 -13304 457 -13266
rect 406 -33184 457 -33146
rect 406 -49727 457 -49689
rect 406 -10180 457 -10142
rect 406 -57395 457 -57357
rect 406 -23457 457 -23419
rect 406 -11742 457 -11704
rect 406 -35527 457 -35489
rect 406 -16357 457 -16319
rect 406 -64850 457 -64812
rect 406 -25729 457 -25691
rect 406 -62436 457 -62398
rect 406 -13517 457 -13479
rect 406 -49656 457 -49618
rect 406 -53845 457 -53807
rect 406 -58176 457 -58138
rect 406 -62365 457 -62327
rect 406 -17280 457 -17242
rect 406 -49585 457 -49547
rect 406 -27291 457 -27253
rect 406 -58886 457 -58848
rect 406 -65986 457 -65948
rect 406 -47313 457 -47275
rect 406 -35740 457 -35702
rect 406 -20333 457 -20295
rect 406 -15718 457 -15680
rect 406 -62862 457 -62824
rect 406 -19055 457 -19017
rect 406 -30060 457 -30022
rect 406 -54271 457 -54233
rect 406 -70885 457 -70847
rect 406 -42272 457 -42234
rect 406 -68542 457 -68504
rect 406 -12594 457 -12556
rect 406 -58744 457 -58706
rect 406 -62507 457 -62469
rect 406 -64353 457 -64315
rect 406 -14440 457 -14402
rect 406 -24877 457 -24839
rect 406 -28853 457 -28815
rect 406 -35385 457 -35347
rect 406 -40852 457 -40814
rect 406 -9683 457 -9645
rect 406 -56330 457 -56292
rect 406 -70956 457 -70918
rect 406 -10464 457 -10426
rect 406 -59738 457 -59700
rect 406 -42414 457 -42376
rect 406 -15292 457 -15254
rect 406 -38651 457 -38613
rect 406 -56046 457 -56008
rect 406 -59028 457 -58990
rect 406 -12736 457 -12698
rect 406 -35314 457 -35276
rect 406 -30841 457 -30803
rect 406 -64282 457 -64244
rect 406 -42556 457 -42518
rect 406 -33397 457 -33359
rect 406 -47455 457 -47417
rect 406 -52283 457 -52245
rect 406 -29563 457 -29525
rect 406 -40142 457 -40104
rect 406 -44615 457 -44577
rect 406 -32971 457 -32933
rect 406 -40355 457 -40317
rect 406 -27646 457 -27608
rect 406 -45112 457 -45074
rect 406 -15576 457 -15538
rect 406 -60590 457 -60552
rect 406 -29776 457 -29738
rect 406 -67619 457 -67581
rect 406 -66696 457 -66658
rect 406 -17564 457 -17526
rect 406 -11032 457 -10994
rect 406 -63146 457 -63108
rect 406 -30912 457 -30874
rect 406 -38438 457 -38400
rect 406 -14511 457 -14473
rect 406 -22605 457 -22567
rect 406 -68471 457 -68433
rect 406 -68968 457 -68930
rect 406 -17990 457 -17952
rect 406 -27504 457 -27466
rect 406 -29989 457 -29951
rect 406 -62720 457 -62682
rect 406 -60377 457 -60339
rect 406 -35598 457 -35560
rect 406 -40284 457 -40246
rect 406 -63856 457 -63818
rect 406 -11103 457 -11065
rect 406 -44970 457 -44932
rect 406 -63288 457 -63250
rect 406 -14866 457 -14828
rect 406 -21469 457 -21431
rect 406 -23599 457 -23561
rect 406 -11884 457 -11846
rect 406 -49017 457 -48979
rect 406 -11529 457 -11491
rect 406 -15434 457 -15396
rect 406 -64069 457 -64031
rect 406 -17209 457 -17171
rect 406 -42698 457 -42660
rect 406 -51715 457 -51677
rect 406 -62649 457 -62611
rect 406 -49230 457 -49192
rect 406 -56117 457 -56079
rect 406 -51644 457 -51606
rect 406 -44473 457 -44435
rect 406 -9825 457 -9787
rect 406 -52141 457 -52103
rect 406 -19126 457 -19088
rect 406 -12807 457 -12769
rect 406 -21185 457 -21147
rect 406 -32261 457 -32223
rect 406 -25019 457 -24981
rect 406 -40781 457 -40743
rect 406 -48946 457 -48908
rect 406 -63643 457 -63605
rect 406 -64637 457 -64599
rect 406 -53916 457 -53878
rect 406 -56543 457 -56505
rect 406 -26936 457 -26898
rect 406 -57466 457 -57428
rect 406 -10677 457 -10639
rect 406 -13588 457 -13550
rect 406 -22747 457 -22709
rect 406 -32190 457 -32152
rect 406 -29847 457 -29809
rect 406 -27717 457 -27679
rect 406 -44899 457 -44861
rect 406 -21398 457 -21360
rect 406 -66767 457 -66729
rect 406 -40497 457 -40459
rect 406 -49088 457 -49050
rect 406 -17422 457 -17384
rect 406 -22534 457 -22496
rect 406 -45183 457 -45145
rect 406 -45467 457 -45429
rect 406 -28640 457 -28602
rect 406 -40426 457 -40388
rect 406 -23741 457 -23703
rect 406 -60306 457 -60268
rect 406 -24593 457 -24555
rect 406 -14937 457 -14899
rect 406 -20475 457 -20437
rect 406 -53774 457 -53736
rect 406 -10890 457 -10852
rect 406 -18132 457 -18094
rect 406 -14724 457 -14686
rect 406 -49301 457 -49263
rect 406 -10748 457 -10710
rect 406 -52212 457 -52174
rect 406 -12239 457 -12201
rect 406 -42201 457 -42163
rect 406 -49798 457 -49760
rect 406 -19268 457 -19230
rect 406 -39929 457 -39891
rect 406 -60519 457 -60481
rect 406 -47526 457 -47488
rect 406 -66199 457 -66161
rect 406 -68258 457 -68220
rect 406 -69891 457 -69853
rect 406 -24735 457 -24697
rect 406 -40071 457 -40033
rect 406 -61371 457 -61333
rect 406 -10393 457 -10355
rect 406 -29705 457 -29667
rect 406 -31835 457 -31797
rect 406 -51289 457 -51251
rect 406 -9470 457 -9432
rect 406 -11671 457 -11633
rect 406 -46958 457 -46920
rect 406 -19197 457 -19159
rect 406 -13943 457 -13905
rect 406 -64495 457 -64457
rect 406 -37586 457 -37548
rect 406 -30770 457 -30732
rect 406 -14298 457 -14260
rect 406 -65773 457 -65735
rect 406 -51502 457 -51464
rect 406 -32048 457 -32010
rect 406 -35669 457 -35631
rect 406 -44544 457 -44506
rect 406 -27078 457 -27040
rect 406 -25871 457 -25833
rect 406 -11955 457 -11917
rect 406 -59596 457 -59558
rect 406 -63217 457 -63179
rect 406 -14014 457 -13976
rect 406 -22676 457 -22638
rect 406 -38509 457 -38471
rect 406 -17848 457 -17810
rect 406 -69039 457 -69001
rect 406 -63927 457 -63889
rect 406 -14369 457 -14331
rect 406 -34249 457 -34211
rect 406 -47171 457 -47133
rect 406 -28427 457 -28389
rect 406 -15150 457 -15112
rect 406 -15221 457 -15183
rect 406 -25800 457 -25762
rect 406 -69749 457 -69711
rect 406 -56401 457 -56363
rect 406 -47100 457 -47062
rect 406 -69252 457 -69214
rect 406 -16712 457 -16674
rect 406 -58318 457 -58280
rect 406 -42840 457 -42802
rect 406 -9328 457 -9290
rect 406 -12026 457 -11988
rect 406 -21114 457 -21076
rect 406 -18984 457 -18946
rect 406 -38012 457 -37974
rect 406 -33042 457 -33004
rect 406 -9541 457 -9503
rect 406 -11387 457 -11349
rect 406 -31196 457 -31158
rect 406 -64566 457 -64528
rect 406 -14227 457 -14189
rect 406 -15505 457 -15467
rect 406 -45041 457 -45003
rect 406 -16286 457 -16248
rect 406 -32332 457 -32294
rect 406 -63501 457 -63463
rect 406 -16925 457 -16887
rect 406 -37799 457 -37761
rect 406 -44402 457 -44364
rect 406 -39858 457 -39820
rect 406 -40639 457 -40601
rect 406 -10251 457 -10213
rect 406 -67548 457 -67510
rect 406 -40213 457 -40175
rect 406 -64708 457 -64670
rect 406 -34178 457 -34140
rect 406 -12878 457 -12840
rect 406 -67051 457 -67013
rect 406 -70672 457 -70634
rect 406 -63714 457 -63676
rect 406 -18061 457 -18023
rect 406 -9754 457 -9716
rect 406 -62223 457 -62185
rect 406 -30699 457 -30661
rect 406 -61158 457 -61120
rect 406 -25942 457 -25904
rect 406 -53703 457 -53665
rect 406 -46674 457 -46636
rect 406 -40923 457 -40885
rect 406 -56614 457 -56576
rect 406 -58247 457 -58209
rect 406 -16428 457 -16390
rect 406 -50011 457 -49973
rect 406 -10109 457 -10071
rect 406 -13233 457 -13195
rect 406 -12452 457 -12414
rect 406 -34604 457 -34566
rect 406 -13446 457 -13408
rect 406 -13375 457 -13337
rect 406 -34320 457 -34282
rect 406 -16641 457 -16603
rect 406 -65915 457 -65877
rect 406 -16570 457 -16532
rect 406 -17493 457 -17455
rect 406 -40000 457 -39962
rect 406 -64779 457 -64741
rect 406 -45396 457 -45358
rect 406 -53561 457 -53523
rect 406 -42130 457 -42092
rect 406 -27575 457 -27537
rect 406 -52070 457 -52032
rect 406 -61087 457 -61049
rect 406 -56188 457 -56150
rect 406 -62294 457 -62256
rect 406 -46887 457 -46849
rect 406 -53987 457 -53949
rect 406 -44686 457 -44648
rect 406 -49514 457 -49476
rect 406 -45325 457 -45287
rect 406 -33468 457 -33430
rect 406 -44828 457 -44790
rect 406 -22321 457 -22283
rect 406 -15789 457 -15751
rect 406 -17067 457 -17029
rect 406 -71098 457 -71060
rect 406 -40568 457 -40530
rect 406 -23670 457 -23632
rect 406 -20404 457 -20366
rect 406 -47668 457 -47630
rect 406 -24948 457 -24910
rect 406 -71169 457 -71131
rect 406 -26155 457 -26117
rect 406 -31125 457 -31087
rect 406 -15079 457 -15041
rect 406 -70814 457 -70776
rect 406 -13730 457 -13692
rect 406 -54058 457 -54020
rect 406 -27362 457 -27324
rect 406 -65844 457 -65806
rect 406 -16215 457 -16177
rect 406 -38154 457 -38116
rect 406 -28782 457 -28744
rect 406 -70104 457 -70066
rect 406 -66128 457 -66090
rect 406 -51857 457 -51819
rect 406 -56472 457 -56434
rect 406 -63430 457 -63392
rect 406 -16073 457 -16035
rect 406 -10322 457 -10284
rect 406 -64921 457 -64883
rect 406 -58815 457 -58777
rect 406 -28498 457 -28460
rect 406 -31054 457 -31016
rect 406 -38296 457 -38258
rect 406 -61229 457 -61191
rect 406 -49372 457 -49334
rect 406 -67690 457 -67652
rect 406 -9612 457 -9574
rect 406 -69181 457 -69143
rect 406 -24522 457 -24484
rect 406 -63785 457 -63747
rect 406 -30983 457 -30945
rect 406 -17777 457 -17739
rect 406 -49940 457 -49902
rect 406 -47739 457 -47701
rect 406 -49159 457 -49121
rect 406 -64211 457 -64173
rect 406 -56259 457 -56221
rect 406 -62791 457 -62753
rect 406 -15860 457 -15822
rect 406 -16783 457 -16745
rect 406 -23386 457 -23348
rect 406 -28924 457 -28886
rect 406 -13872 457 -13834
rect 406 -17138 457 -17100
rect 406 -9896 457 -9858
rect 406 -24664 457 -24626
rect 406 -12310 457 -12272
rect 406 -66057 457 -66019
rect 406 -27220 457 -27182
rect 406 -16499 457 -16461
rect 406 -70033 457 -69995
rect 406 -46745 457 -46707
rect 406 -66838 457 -66800
rect 406 -47242 457 -47204
rect 406 -17706 457 -17668
rect 406 -12949 457 -12911
rect 406 -66909 457 -66871
rect 406 -37657 457 -37619
rect 406 -34107 457 -34069
rect 406 -13020 457 -12982
rect 406 -9115 457 -9077
rect 406 -16854 457 -16816
rect 406 -51431 457 -51393
rect 406 -9186 457 -9148
rect 406 -64992 457 -64954
rect 406 -26084 457 -26046
rect 406 -33255 457 -33217
rect 406 -71027 457 -70989
rect 406 -21540 457 -21502
rect 406 -33113 457 -33075
rect 406 -62578 457 -62540
rect 406 -11600 457 -11562
rect 406 -38367 457 -38329
rect 406 -18913 457 -18875
rect 406 -67761 457 -67723
rect 406 -20049 457 -20011
rect 406 -64140 457 -64102
rect 406 -14653 457 -14615
rect 406 -63998 457 -63960
rect 406 -22250 457 -22212
rect 406 -10606 457 -10568
rect 406 -21327 457 -21289
rect 406 -20262 457 -20224
rect 406 -12381 457 -12343
rect 406 -18842 457 -18804
rect 406 -11174 457 -11136
rect 406 -17919 457 -17881
rect 406 -10961 457 -10923
rect 406 -14085 457 -14047
rect 406 -63359 457 -63321
rect 406 -69110 457 -69072
rect 406 -69820 457 -69782
rect 406 -40710 457 -40672
rect 406 -42982 457 -42944
rect 406 -15931 457 -15893
rect 406 -23812 457 -23774
rect 406 -21256 457 -21218
rect 406 -22392 457 -22354
rect 406 -32119 457 -32081
rect 406 -45254 457 -45216
rect 406 -65063 457 -65025
rect 406 -14156 457 -14118
rect 406 -12665 457 -12627
rect 406 -11813 457 -11775
rect 406 -67477 457 -67439
rect 406 -13091 457 -13053
rect 406 -68329 457 -68291
rect 406 -68400 457 -68362
rect 406 -35456 457 -35418
rect 406 -35243 457 -35205
rect 406 -31906 457 -31868
rect 406 -54129 457 -54091
rect 406 -49443 457 -49405
rect 406 -23528 457 -23490
rect 406 -11458 457 -11420
rect 406 -27149 457 -27111
rect 406 -17351 457 -17313
rect 406 -71240 457 -71202
rect 406 -61300 457 -61262
rect 406 -47029 457 -46991
rect 406 -37870 457 -37832
rect 406 -28569 457 -28531
rect 406 -69962 457 -69924
rect 406 -58105 457 -58067
rect 406 -63004 457 -62966
rect 406 -19978 457 -19940
rect 406 -34462 457 -34424
rect 406 -27433 457 -27395
rect 406 -54342 457 -54304
rect 406 -23883 457 -23845
rect 406 -12097 457 -12059
rect 406 -20120 457 -20082
rect 406 -14795 457 -14757
rect 406 -49869 457 -49831
rect 406 -63075 457 -63037
rect 406 -11316 457 -11278
rect 406 -34533 457 -34495
rect 406 -27007 457 -26969
rect 406 -61513 457 -61475
rect 406 -25658 457 -25620
rect 406 -59525 457 -59487
rect 406 -33326 457 -33288
rect 406 -46816 457 -46778
rect 406 -61442 457 -61404
rect 406 -15647 457 -15609
rect 406 -59667 457 -59629
rect 406 -29918 457 -29880
rect 406 -57253 457 -57215
rect 406 -13659 457 -13621
rect 406 -9967 457 -9929
rect 406 -54413 457 -54375
rect 406 -47597 457 -47559
rect 406 -57537 457 -57499
rect 406 -57324 457 -57286
rect 406 -58034 457 -57996
rect 406 -10038 457 -10000
rect 406 -60235 457 -60197
rect 406 -13162 457 -13124
rect 406 -26865 457 -26827
rect 406 -64424 457 -64386
rect 406 -16002 457 -15964
rect 406 -47384 457 -47346
rect 406 -38083 457 -38045
rect 406 -9399 457 -9361
rect 406 -51573 457 -51535
rect 406 -16996 457 -16958
rect 406 -51928 457 -51890
rect 406 -12523 457 -12485
rect 406 -20191 457 -20153
rect 406 -38225 457 -38187
rect 406 -21611 457 -21573
rect 406 -28711 457 -28673
rect 406 -26794 457 -26756
rect 406 -38580 457 -38542
rect 406 -37728 457 -37690
rect 406 -17635 457 -17597
rect 406 -59809 457 -59771
rect 406 -34391 457 -34353
rect 406 -13801 457 -13763
rect 406 -60448 457 -60410
rect 406 -42343 457 -42305
rect 406 -53632 457 -53594
rect 406 -12168 457 -12130
rect 406 -14582 457 -14544
rect 406 -51999 457 -51961
rect 406 -42485 457 -42447
rect 406 -54484 457 -54446
rect 406 -51786 457 -51748
rect 406 -63572 457 -63534
rect 406 -44757 457 -44719
rect 406 -42769 457 -42731
rect 406 -19339 457 -19301
rect 240 -29634 291 -29596
rect 240 -10535 291 -10497
rect 240 -66980 291 -66942
rect 240 -15363 291 -15325
rect 240 -34675 291 -34637
rect 240 -53490 291 -53452
rect 240 -54200 291 -54162
rect 240 -57182 291 -57144
rect 240 -30628 291 -30590
rect 240 -11245 291 -11207
rect 240 -28143 291 -28105
rect 240 -39432 291 -39394
rect 240 -56827 291 -56789
rect 240 -31977 291 -31939
rect 240 -27788 291 -27750
rect 240 -15008 291 -14970
rect 240 -48520 291 -48482
rect 240 -68684 291 -68646
rect 240 -16144 291 -16106
rect 240 -10819 291 -10781
rect 240 -59951 291 -59913
rect 240 -65347 291 -65309
rect 240 -24806 291 -24768
rect 240 -22463 291 -22425
rect 240 -9257 291 -9219
rect 240 -62933 291 -62895
rect 240 -58957 291 -58919
rect 240 -13304 291 -13266
rect 240 -24451 291 -24413
rect 240 -43692 291 -43654
rect 240 -49727 291 -49689
rect 240 -10180 291 -10142
rect 240 -57395 291 -57357
rect 240 -11742 291 -11704
rect 240 -16357 291 -16319
rect 240 -64850 291 -64812
rect 240 -24025 291 -23987
rect 240 -58602 291 -58564
rect 240 -62436 291 -62398
rect 240 -13517 291 -13479
rect 240 -49656 291 -49618
rect 240 -53845 291 -53807
rect 240 -62365 291 -62327
rect 240 -17280 291 -17242
rect 240 -70388 291 -70350
rect 240 -49585 291 -49547
rect 240 -43479 291 -43441
rect 240 -22037 291 -21999
rect 240 -27291 291 -27253
rect 240 -58886 291 -58848
rect 240 -38935 291 -38897
rect 240 -28072 291 -28034
rect 240 -52780 291 -52742
rect 240 -20333 291 -20295
rect 240 -15718 291 -15680
rect 240 -62862 291 -62824
rect 240 -52567 291 -52529
rect 240 -43408 291 -43370
rect 240 -30060 291 -30022
rect 240 -54271 291 -54233
rect 240 -61939 291 -61901
rect 240 -35172 291 -35134
rect 240 -67406 291 -67368
rect 240 -43905 291 -43867
rect 240 -68542 291 -68504
rect 240 -12594 291 -12556
rect 240 -26297 291 -26259
rect 240 -58744 291 -58706
rect 240 -62507 291 -62469
rect 240 -19694 291 -19656
rect 240 -64353 291 -64315
rect 240 -14440 291 -14402
rect 240 -24877 291 -24839
rect 240 -27930 291 -27892
rect 240 -40852 291 -40814
rect 240 -9683 291 -9645
rect 240 -10464 291 -10426
rect 240 -15292 291 -15254
rect 240 -59028 291 -58990
rect 240 -12736 291 -12698
rect 240 -34746 291 -34708
rect 240 -26510 291 -26472
rect 240 -34959 291 -34921
rect 240 -64282 291 -64244
rect 240 -29563 291 -29525
rect 240 -40142 291 -40104
rect 240 -48733 291 -48695
rect 240 -44615 291 -44577
rect 240 -40355 291 -40317
rect 240 -27646 291 -27608
rect 240 -45112 291 -45074
rect 240 -15576 291 -15538
rect 240 -60590 291 -60552
rect 240 -68755 291 -68717
rect 240 -29776 291 -29738
rect 240 -32758 291 -32720
rect 240 -39645 291 -39607
rect 240 -32687 291 -32649
rect 240 -66696 291 -66658
rect 240 -21753 291 -21715
rect 240 -17564 291 -17526
rect 240 -65276 291 -65238
rect 240 -11032 291 -10994
rect 240 -63146 291 -63108
rect 240 -58531 291 -58493
rect 240 -53064 291 -53026
rect 240 -14511 291 -14473
rect 240 -22605 291 -22567
rect 240 -21966 291 -21928
rect 240 -68471 291 -68433
rect 240 -65631 291 -65593
rect 240 -17990 291 -17952
rect 240 -27504 291 -27466
rect 240 -29989 291 -29951
rect 240 -32474 291 -32436
rect 240 -62720 291 -62682
rect 240 -60377 291 -60339
rect 240 -63856 291 -63818
rect 240 -40284 291 -40246
rect 240 -11103 291 -11065
rect 240 -44970 291 -44932
rect 240 -63288 291 -63250
rect 240 -14866 291 -14828
rect 240 -62081 291 -62043
rect 240 -11884 291 -11846
rect 240 -49017 291 -48979
rect 240 -11529 291 -11491
rect 240 -15434 291 -15396
rect 240 -64069 291 -64031
rect 240 -32403 291 -32365
rect 240 -17209 291 -17171
rect 240 -47881 291 -47843
rect 240 -48449 291 -48411
rect 240 -62649 291 -62611
rect 240 -49230 291 -49192
rect 240 -68613 291 -68575
rect 240 -44473 291 -44435
rect 240 -9825 291 -9787
rect 240 -52638 291 -52600
rect 240 -70459 291 -70421
rect 240 -12807 291 -12769
rect 240 -32261 291 -32223
rect 240 -44189 291 -44151
rect 240 -57040 291 -57002
rect 240 -25019 291 -24981
rect 240 -40781 291 -40743
rect 240 -48946 291 -48908
rect 240 -63643 291 -63605
rect 240 -64637 291 -64599
rect 240 -53916 291 -53878
rect 240 -39077 291 -39039
rect 240 -19907 291 -19869
rect 240 -26936 291 -26898
rect 240 -57466 291 -57428
rect 240 -10677 291 -10639
rect 240 -65205 291 -65167
rect 240 -13588 291 -13550
rect 240 -22747 291 -22709
rect 240 -32190 291 -32152
rect 240 -29847 291 -29809
rect 240 -48023 291 -47985
rect 240 -27717 291 -27679
rect 240 -62010 291 -61972
rect 240 -44899 291 -44861
rect 240 -66767 291 -66729
rect 240 -58389 291 -58351
rect 240 -40497 291 -40459
rect 240 -49088 291 -49050
rect 240 -17422 291 -17384
rect 240 -24096 291 -24058
rect 240 -47952 291 -47914
rect 240 -30131 291 -30093
rect 240 -22534 291 -22496
rect 240 -45183 291 -45145
rect 240 -45467 291 -45429
rect 240 -60164 291 -60126
rect 240 -40426 291 -40388
rect 240 -60306 291 -60268
rect 240 -24593 291 -24555
rect 240 -14937 291 -14899
rect 240 -32545 291 -32507
rect 240 -20475 291 -20437
rect 240 -21682 291 -21644
rect 240 -53774 291 -53736
rect 240 -10890 291 -10852
rect 240 -18132 291 -18094
rect 240 -14724 291 -14686
rect 240 -49301 291 -49263
rect 240 -10748 291 -10710
rect 240 -12239 291 -12201
rect 240 -24380 291 -24342
rect 240 -49798 291 -49760
rect 240 -39929 291 -39891
rect 240 -19410 291 -19372
rect 240 -60519 291 -60481
rect 240 -68258 291 -68220
rect 240 -22179 291 -22141
rect 240 -69891 291 -69853
rect 240 -24735 291 -24697
rect 240 -39503 291 -39465
rect 240 -19481 291 -19443
rect 240 -40071 291 -40033
rect 240 -26652 291 -26614
rect 240 -56685 291 -56647
rect 240 -10393 291 -10355
rect 240 -26368 291 -26330
rect 240 -29705 291 -29667
rect 240 -31835 291 -31797
rect 240 -9470 291 -9432
rect 240 -11671 291 -11633
rect 240 -60093 291 -60055
rect 240 -48165 291 -48127
rect 240 -64495 291 -64457
rect 240 -13943 291 -13905
rect 240 -53419 291 -53381
rect 240 -14298 291 -14260
rect 240 -32048 291 -32010
rect 240 -44544 291 -44506
rect 240 -27078 291 -27040
rect 240 -59880 291 -59842
rect 240 -24167 291 -24129
rect 240 -39290 291 -39252
rect 240 -11955 291 -11917
rect 240 -63217 291 -63179
rect 240 -14014 291 -13976
rect 240 -22676 291 -22638
rect 240 -17848 291 -17810
rect 240 -35030 291 -34992
rect 240 -56898 291 -56860
rect 240 -60022 291 -59984
rect 240 -63927 291 -63889
rect 240 -14369 291 -14331
rect 240 -34249 291 -34211
rect 240 -24309 291 -24271
rect 240 -15150 291 -15112
rect 240 -15221 291 -15183
rect 240 -70530 291 -70492
rect 240 -69749 291 -69711
rect 240 -52496 291 -52458
rect 240 -44260 291 -44222
rect 240 -16712 291 -16674
rect 240 -9328 291 -9290
rect 240 -12026 291 -11988
rect 240 -52922 291 -52884
rect 240 -9541 291 -9503
rect 240 -11387 291 -11349
rect 240 -64566 291 -64528
rect 240 -14227 291 -14189
rect 240 -24238 291 -24200
rect 240 -26581 291 -26543
rect 240 -15505 291 -15467
rect 240 -45041 291 -45003
rect 240 -65418 291 -65380
rect 240 -16286 291 -16248
rect 240 -32332 291 -32294
rect 240 -63501 291 -63463
rect 240 -26723 291 -26685
rect 240 -16925 291 -16887
rect 240 -48591 291 -48553
rect 240 -44402 291 -44364
rect 240 -68897 291 -68859
rect 240 -39858 291 -39820
rect 240 -40639 291 -40601
rect 240 -10251 291 -10213
rect 240 -40213 291 -40175
rect 240 -64708 291 -64670
rect 240 -34178 291 -34140
rect 240 -12878 291 -12840
rect 240 -47810 291 -47772
rect 240 -67051 291 -67013
rect 240 -63714 291 -63676
rect 240 -18061 291 -18023
rect 240 -9754 291 -9716
rect 240 -21824 291 -21786
rect 240 -62223 291 -62185
rect 240 -53703 291 -53665
rect 240 -40923 291 -40885
rect 240 -70317 291 -70279
rect 240 -16428 291 -16390
rect 240 -35101 291 -35063
rect 240 -50011 291 -49973
rect 240 -10109 291 -10071
rect 240 -13233 291 -13195
rect 240 -12452 291 -12414
rect 240 -34604 291 -34566
rect 240 -13446 291 -13408
rect 240 -13375 291 -13337
rect 240 -34320 291 -34282
rect 240 -16641 291 -16603
rect 240 -16570 291 -16532
rect 240 -17493 291 -17455
rect 240 -40000 291 -39962
rect 240 -48378 291 -48340
rect 240 -64779 291 -64741
rect 240 -45396 291 -45358
rect 240 -38864 291 -38826
rect 240 -53561 291 -53523
rect 240 -27575 291 -27537
rect 240 -62294 291 -62256
rect 240 -68826 291 -68788
rect 240 -39006 291 -38968
rect 240 -48236 291 -48198
rect 240 -53987 291 -53949
rect 240 -58460 291 -58422
rect 240 -44686 291 -44648
rect 240 -32900 291 -32862
rect 240 -49514 291 -49476
rect 240 -30486 291 -30448
rect 240 -45325 291 -45287
rect 240 -44828 291 -44790
rect 240 -22321 291 -22283
rect 240 -15789 291 -15751
rect 240 -17067 291 -17029
rect 240 -40568 291 -40530
rect 240 -52851 291 -52813
rect 240 -30344 291 -30306
rect 240 -20404 291 -20366
rect 240 -70246 291 -70208
rect 240 -24948 291 -24910
rect 240 -28214 291 -28176
rect 240 -53206 291 -53168
rect 240 -32616 291 -32578
rect 240 -27859 291 -27821
rect 240 -15079 291 -15041
rect 240 -13730 291 -13692
rect 240 -54058 291 -54020
rect 240 -61868 291 -61830
rect 240 -70601 291 -70563
rect 240 -27362 291 -27324
rect 240 -61726 291 -61688
rect 240 -39361 291 -39323
rect 240 -16215 291 -16177
rect 240 -19552 291 -19514
rect 240 -39219 291 -39181
rect 240 -19623 291 -19585
rect 240 -70104 291 -70066
rect 240 -63430 291 -63392
rect 240 -16073 291 -16035
rect 240 -10322 291 -10284
rect 240 -64921 291 -64883
rect 240 -58815 291 -58777
rect 240 -43976 291 -43938
rect 240 -65134 291 -65096
rect 240 -67335 291 -67297
rect 240 -48804 291 -48766
rect 240 -57111 291 -57073
rect 240 -26226 291 -26188
rect 240 -49372 291 -49334
rect 240 -21895 291 -21857
rect 240 -9612 291 -9574
rect 240 -67122 291 -67084
rect 240 -61797 291 -61759
rect 240 -24522 291 -24484
rect 240 -63785 291 -63747
rect 240 -17777 291 -17739
rect 240 -52425 291 -52387
rect 240 -22108 291 -22070
rect 240 -53348 291 -53310
rect 240 -43266 291 -43228
rect 240 -49940 291 -49902
rect 240 -49159 291 -49121
rect 240 -64211 291 -64173
rect 240 -62791 291 -62753
rect 240 -15860 291 -15822
rect 240 -16783 291 -16745
rect 240 -13872 291 -13834
rect 240 -17138 291 -17100
rect 240 -9896 291 -9858
rect 240 -24664 291 -24626
rect 240 -39574 291 -39536
rect 240 -12310 291 -12272
rect 240 -34817 291 -34779
rect 240 -27220 291 -27182
rect 240 -16499 291 -16461
rect 240 -70033 291 -69995
rect 240 -66838 291 -66800
rect 240 -28285 291 -28247
rect 240 -19836 291 -19798
rect 240 -44118 291 -44080
rect 240 -17706 291 -17668
rect 240 -12949 291 -12911
rect 240 -66909 291 -66871
rect 240 -34107 291 -34069
rect 240 -13020 291 -12982
rect 240 -53277 291 -53239
rect 240 -9115 291 -9077
rect 240 -16854 291 -16816
rect 240 -9186 291 -9148
rect 240 -64992 291 -64954
rect 240 -53135 291 -53097
rect 240 -70175 291 -70137
rect 240 -30202 291 -30164
rect 240 -62578 291 -62540
rect 240 -11600 291 -11562
rect 240 -20049 291 -20011
rect 240 -38793 291 -38755
rect 240 -64140 291 -64102
rect 240 -14653 291 -14615
rect 240 -63998 291 -63960
rect 240 -22250 291 -22212
rect 240 -10606 291 -10568
rect 240 -20262 291 -20224
rect 240 -12381 291 -12343
rect 240 -11174 291 -11136
rect 240 -17919 291 -17881
rect 240 -10961 291 -10923
rect 240 -14085 291 -14047
rect 240 -63359 291 -63321
rect 240 -39148 291 -39110
rect 240 -69820 291 -69782
rect 240 -40710 291 -40672
rect 240 -15931 291 -15893
rect 240 -61584 291 -61546
rect 240 -67264 291 -67226
rect 240 -62152 291 -62114
rect 240 -30557 291 -30519
rect 240 -22392 291 -22354
rect 240 -32119 291 -32081
rect 240 -45254 291 -45216
rect 240 -48094 291 -48056
rect 240 -65063 291 -65025
rect 240 -14156 291 -14118
rect 240 -39787 291 -39749
rect 240 -12665 291 -12627
rect 240 -11813 291 -11775
rect 240 -34888 291 -34850
rect 240 -48307 291 -48269
rect 240 -13091 291 -13053
rect 240 -68329 291 -68291
rect 240 -68400 291 -68362
rect 240 -48662 291 -48624
rect 240 -30273 291 -30235
rect 240 -38722 291 -38684
rect 240 -43621 291 -43583
rect 240 -52709 291 -52671
rect 240 -31906 291 -31868
rect 240 -54129 291 -54091
rect 240 -43337 291 -43299
rect 240 -49443 291 -49405
rect 240 -58673 291 -58635
rect 240 -43763 291 -43725
rect 240 -11458 291 -11420
rect 240 -27149 291 -27111
rect 240 -17351 291 -17313
rect 240 -43550 291 -43512
rect 240 -69962 291 -69924
rect 240 -28356 291 -28318
rect 240 -63004 291 -62966
rect 240 -19978 291 -19940
rect 240 -34462 291 -34424
rect 240 -26439 291 -26401
rect 240 -56969 291 -56931
rect 240 -27433 291 -27395
rect 240 -65560 291 -65522
rect 240 -54342 291 -54304
rect 240 -12097 291 -12059
rect 240 -20120 291 -20082
rect 240 -14795 291 -14757
rect 240 -49869 291 -49831
rect 240 -63075 291 -63037
rect 240 -28001 291 -27963
rect 240 -11316 291 -11278
rect 240 -34533 291 -34495
rect 240 -61655 291 -61617
rect 240 -27007 291 -26969
rect 240 -15647 291 -15609
rect 240 -29918 291 -29880
rect 240 -48875 291 -48837
rect 240 -43834 291 -43796
rect 240 -57253 291 -57215
rect 240 -65702 291 -65664
rect 240 -13659 291 -13621
rect 240 -9967 291 -9929
rect 240 -54413 291 -54375
rect 240 -52354 291 -52316
rect 240 -57537 291 -57499
rect 240 -57324 291 -57286
rect 240 -32829 291 -32791
rect 240 -10038 291 -10000
rect 240 -30415 291 -30377
rect 240 -60235 291 -60197
rect 240 -13162 291 -13124
rect 240 -26865 291 -26827
rect 240 -64424 291 -64386
rect 240 -16002 291 -15964
rect 240 -9399 291 -9361
rect 240 -16996 291 -16958
rect 240 -12523 291 -12485
rect 240 -20191 291 -20153
rect 240 -26794 291 -26756
rect 240 -44331 291 -44293
rect 240 -44047 291 -44009
rect 240 -23954 291 -23916
rect 240 -17635 291 -17597
rect 240 -65489 291 -65451
rect 240 -34391 291 -34353
rect 240 -13801 291 -13763
rect 240 -60448 291 -60410
rect 240 -53632 291 -53594
rect 240 -12168 291 -12130
rect 240 -14582 291 -14544
rect 240 -39716 291 -39678
rect 240 -67193 291 -67155
rect 240 -19765 291 -19727
rect 240 -54484 291 -54446
rect 240 -63572 291 -63534
rect 240 -44757 291 -44719
rect 240 -52993 291 -52955
rect 240 -56756 291 -56718
rect 157 -29208 208 -29170
rect 157 -42911 208 -42873
rect 157 -10535 208 -10497
rect 157 -51360 208 -51322
rect 157 -42627 208 -42589
rect 157 -15363 208 -15325
rect 157 -26013 208 -25975
rect 157 -53490 208 -53452
rect 157 -41633 208 -41595
rect 157 -20901 208 -20863
rect 157 -54200 208 -54162
rect 157 -43053 208 -43015
rect 157 -11245 208 -11207
rect 157 -41349 208 -41311
rect 157 -28143 208 -28105
rect 157 -31977 208 -31939
rect 157 -41420 208 -41382
rect 157 -43124 208 -43086
rect 157 -27788 208 -27750
rect 157 -15008 208 -14970
rect 157 -68684 208 -68646
rect 157 -16144 208 -16106
rect 157 -10819 208 -10781
rect 157 -65347 208 -65309
rect 157 -43195 208 -43157
rect 157 -51218 208 -51180
rect 157 -22463 208 -22425
rect 157 -9257 208 -9219
rect 157 -62933 208 -62895
rect 157 -58957 208 -58919
rect 157 -13304 208 -13266
rect 157 -33184 208 -33146
rect 157 -20688 208 -20650
rect 157 -40994 208 -40956
rect 157 -43692 208 -43654
rect 157 -10180 208 -10142
rect 157 -29350 208 -29312
rect 157 -25374 208 -25336
rect 157 -11742 208 -11704
rect 157 -16357 208 -16319
rect 157 -64850 208 -64812
rect 157 -25729 208 -25691
rect 157 -58602 208 -58564
rect 157 -20759 208 -20721
rect 157 -62436 208 -62398
rect 157 -66341 208 -66303
rect 157 -13517 208 -13479
rect 157 -53845 208 -53807
rect 157 -58176 208 -58138
rect 157 -62365 208 -62327
rect 157 -17280 208 -17242
rect 157 -51076 208 -51038
rect 157 -43479 208 -43441
rect 157 -22037 208 -21999
rect 157 -27291 208 -27253
rect 157 -58886 208 -58848
rect 157 -65986 208 -65948
rect 157 -52780 208 -52742
rect 157 -28072 208 -28034
rect 157 -51005 208 -50967
rect 157 -15718 208 -15680
rect 157 -62862 208 -62824
rect 157 -52567 208 -52529
rect 157 -43408 208 -43370
rect 157 -54271 208 -54233
rect 157 -61939 208 -61901
rect 157 -50579 208 -50541
rect 157 -43905 208 -43867
rect 157 -42272 208 -42234
rect 157 -50934 208 -50896
rect 157 -68542 208 -68504
rect 157 -12594 208 -12556
rect 157 -26297 208 -26259
rect 157 -58744 208 -58706
rect 157 -62507 208 -62469
rect 157 -64353 208 -64315
rect 157 -14440 208 -14402
rect 157 -66483 208 -66445
rect 157 -27930 208 -27892
rect 157 -28853 208 -28815
rect 157 -9683 208 -9645
rect 157 -10464 208 -10426
rect 157 -20546 208 -20508
rect 157 -50863 208 -50825
rect 157 -42414 208 -42376
rect 157 -60874 208 -60836
rect 157 -15292 208 -15254
rect 157 -41278 208 -41240
rect 157 -41065 208 -41027
rect 157 -59028 208 -58990
rect 157 -12736 208 -12698
rect 157 -25516 208 -25478
rect 157 -26510 208 -26472
rect 157 -60803 208 -60765
rect 157 -64282 208 -64244
rect 157 -42556 208 -42518
rect 157 -33397 208 -33359
rect 157 -52283 208 -52245
rect 157 -69394 208 -69356
rect 157 -44615 208 -44577
rect 157 -32971 208 -32933
rect 157 -27646 208 -27608
rect 157 -45112 208 -45074
rect 157 -15576 208 -15538
rect 157 -41917 208 -41879
rect 157 -68755 208 -68717
rect 157 -32758 208 -32720
rect 157 -50721 208 -50683
rect 157 -32687 208 -32649
rect 157 -21753 208 -21715
rect 157 -17564 208 -17526
rect 157 -65276 208 -65238
rect 157 -11032 208 -10994
rect 157 -63146 208 -63108
rect 157 -50153 208 -50115
rect 157 -58531 208 -58493
rect 157 -53064 208 -53026
rect 157 -14511 208 -14473
rect 157 -22605 208 -22567
rect 157 -21966 208 -21928
rect 157 -68471 208 -68433
rect 157 -65631 208 -65593
rect 157 -68968 208 -68930
rect 157 -17990 208 -17952
rect 157 -27504 208 -27466
rect 157 -32474 208 -32436
rect 157 -62720 208 -62682
rect 157 -63856 208 -63818
rect 157 -11103 208 -11065
rect 157 -44970 208 -44932
rect 157 -63288 208 -63250
rect 157 -14866 208 -14828
rect 157 -21469 208 -21431
rect 157 -62081 208 -62043
rect 157 -11884 208 -11846
rect 157 -11529 208 -11491
rect 157 -15434 208 -15396
rect 157 -64069 208 -64031
rect 157 -32403 208 -32365
rect 157 -17209 208 -17171
rect 157 -42698 208 -42660
rect 157 -51715 208 -51677
rect 157 -33894 208 -33856
rect 157 -62649 208 -62611
rect 157 -25587 208 -25549
rect 157 -68613 208 -68575
rect 157 -51644 208 -51606
rect 157 -44473 208 -44435
rect 157 -9825 208 -9787
rect 157 -52141 208 -52103
rect 157 -52638 208 -52600
rect 157 -12807 208 -12769
rect 157 -21185 208 -21147
rect 157 -32261 208 -32223
rect 157 -44189 208 -44151
rect 157 -33539 208 -33501
rect 157 -63643 208 -63605
rect 157 -64637 208 -64599
rect 157 -25232 208 -25194
rect 157 -53916 208 -53878
rect 157 -26936 208 -26898
rect 157 -33681 208 -33643
rect 157 -10677 208 -10639
rect 157 -65205 208 -65167
rect 157 -13588 208 -13550
rect 157 -22747 208 -22709
rect 157 -32190 208 -32152
rect 157 -27717 208 -27679
rect 157 -50437 208 -50399
rect 157 -62010 208 -61972
rect 157 -44899 208 -44861
rect 157 -21398 208 -21360
rect 157 -58389 208 -58351
rect 157 -17422 208 -17384
rect 157 -22534 208 -22496
rect 157 -45183 208 -45145
rect 157 -45467 208 -45429
rect 157 -28640 208 -28602
rect 157 -29066 208 -29028
rect 157 -14937 208 -14899
rect 157 -32545 208 -32507
rect 157 -21682 208 -21644
rect 157 -53774 208 -53736
rect 157 -10890 208 -10852
rect 157 -18132 208 -18094
rect 157 -14724 208 -14686
rect 157 -10748 208 -10710
rect 157 -33610 208 -33572
rect 157 -52212 208 -52174
rect 157 -12239 208 -12201
rect 157 -33965 208 -33927
rect 157 -41775 208 -41737
rect 157 -42201 208 -42163
rect 157 -50508 208 -50470
rect 157 -33823 208 -33785
rect 157 -41491 208 -41453
rect 157 -25090 208 -25052
rect 157 -68258 208 -68220
rect 157 -66199 208 -66161
rect 157 -22179 208 -22141
rect 157 -26652 208 -26614
rect 157 -21043 208 -21005
rect 157 -61371 208 -61333
rect 157 -10393 208 -10355
rect 157 -26368 208 -26330
rect 157 -31835 208 -31797
rect 157 -51289 208 -51251
rect 157 -29279 208 -29241
rect 157 -9470 208 -9432
rect 157 -11671 208 -11633
rect 157 -64495 208 -64457
rect 157 -13943 208 -13905
rect 157 -53419 208 -53381
rect 157 -14298 208 -14260
rect 157 -65773 208 -65735
rect 157 -51502 208 -51464
rect 157 -32048 208 -32010
rect 157 -44544 208 -44506
rect 157 -27078 208 -27040
rect 157 -25871 208 -25833
rect 157 -29137 208 -29099
rect 157 -11955 208 -11917
rect 157 -61016 208 -60978
rect 157 -50650 208 -50612
rect 157 -63217 208 -63179
rect 157 -14014 208 -13976
rect 157 -22676 208 -22638
rect 157 -17848 208 -17810
rect 157 -41136 208 -41098
rect 157 -60732 208 -60694
rect 157 -69039 208 -69001
rect 157 -63927 208 -63889
rect 157 -14369 208 -14331
rect 157 -28427 208 -28389
rect 157 -15150 208 -15112
rect 157 -15221 208 -15183
rect 157 -25800 208 -25762
rect 157 -52496 208 -52458
rect 157 -57608 208 -57570
rect 157 -44260 208 -44222
rect 157 -69252 208 -69214
rect 157 -16712 208 -16674
rect 157 -58318 208 -58280
rect 157 -42840 208 -42802
rect 157 -50295 208 -50257
rect 157 -9328 208 -9290
rect 157 -12026 208 -11988
rect 157 -21114 208 -21076
rect 157 -52922 208 -52884
rect 157 -33042 208 -33004
rect 157 -9541 208 -9503
rect 157 -11387 208 -11349
rect 157 -64566 208 -64528
rect 157 -14227 208 -14189
rect 157 -26581 208 -26543
rect 157 -15505 208 -15467
rect 157 -45041 208 -45003
rect 157 -65418 208 -65380
rect 157 -16286 208 -16248
rect 157 -32332 208 -32294
rect 157 -60661 208 -60623
rect 157 -63501 208 -63463
rect 157 -26723 208 -26685
rect 157 -16925 208 -16887
rect 157 -41207 208 -41169
rect 157 -44402 208 -44364
rect 157 -68897 208 -68859
rect 157 -10251 208 -10213
rect 157 -60945 208 -60907
rect 157 -64708 208 -64670
rect 157 -12878 208 -12840
rect 157 -63714 208 -63676
rect 157 -18061 208 -18023
rect 157 -9754 208 -9716
rect 157 -21824 208 -21786
rect 157 -62223 208 -62185
rect 157 -61158 208 -61120
rect 157 -25942 208 -25904
rect 157 -53703 208 -53665
rect 157 -58247 208 -58209
rect 157 -16428 208 -16390
rect 157 -10109 208 -10071
rect 157 -13233 208 -13195
rect 157 -12452 208 -12414
rect 157 -13446 208 -13408
rect 157 -50224 208 -50186
rect 157 -57679 208 -57641
rect 157 -13375 208 -13337
rect 157 -65915 208 -65877
rect 157 -16641 208 -16603
rect 157 -50792 208 -50754
rect 157 -16570 208 -16532
rect 157 -17493 208 -17455
rect 157 -64779 208 -64741
rect 157 -45396 208 -45358
rect 157 -53561 208 -53523
rect 157 -42130 208 -42092
rect 157 -27575 208 -27537
rect 157 -29421 208 -29383
rect 157 -52070 208 -52032
rect 157 -61087 208 -61049
rect 157 -62294 208 -62256
rect 157 -68826 208 -68788
rect 157 -53987 208 -53949
rect 157 -57963 208 -57925
rect 157 -58460 208 -58422
rect 157 -44686 208 -44648
rect 157 -32900 208 -32862
rect 157 -45325 208 -45287
rect 157 -33468 208 -33430
rect 157 -44828 208 -44790
rect 157 -22321 208 -22283
rect 157 -15789 208 -15751
rect 157 -17067 208 -17029
rect 157 -28995 208 -28957
rect 157 -52851 208 -52813
rect 157 -69323 208 -69285
rect 157 -26155 208 -26117
rect 157 -28214 208 -28176
rect 157 -53206 208 -53168
rect 157 -32616 208 -32578
rect 157 -27859 208 -27821
rect 157 -15079 208 -15041
rect 157 -25303 208 -25265
rect 157 -13730 208 -13692
rect 157 -54058 208 -54020
rect 157 -61868 208 -61830
rect 157 -27362 208 -27324
rect 157 -61726 208 -61688
rect 157 -65844 208 -65806
rect 157 -16215 208 -16177
rect 157 -41846 208 -41808
rect 157 -25445 208 -25407
rect 157 -57821 208 -57783
rect 157 -28782 208 -28744
rect 157 -66128 208 -66090
rect 157 -51857 208 -51819
rect 157 -63430 208 -63392
rect 157 -16073 208 -16035
rect 157 -10322 208 -10284
rect 157 -41988 208 -41950
rect 157 -64921 208 -64883
rect 157 -58815 208 -58777
rect 157 -28498 208 -28460
rect 157 -43976 208 -43938
rect 157 -65134 208 -65096
rect 157 -26226 208 -26188
rect 157 -61229 208 -61191
rect 157 -21895 208 -21857
rect 157 -57750 208 -57712
rect 157 -9612 208 -9574
rect 157 -69181 208 -69143
rect 157 -61797 208 -61759
rect 157 -63785 208 -63747
rect 157 -17777 208 -17739
rect 157 -52425 208 -52387
rect 157 -22108 208 -22070
rect 157 -53348 208 -53310
rect 157 -43266 208 -43228
rect 157 -25161 208 -25123
rect 157 -64211 208 -64173
rect 157 -62791 208 -62753
rect 157 -15860 208 -15822
rect 157 -16783 208 -16745
rect 157 -28924 208 -28886
rect 157 -13872 208 -13834
rect 157 -17138 208 -17100
rect 157 -9896 208 -9858
rect 157 -12310 208 -12272
rect 157 -66057 208 -66019
rect 157 -27220 208 -27182
rect 157 -16499 208 -16461
rect 157 -34036 208 -33998
rect 157 -28285 208 -28247
rect 157 -44118 208 -44080
rect 157 -17706 208 -17668
rect 157 -12949 208 -12911
rect 157 -41562 208 -41524
rect 157 -13020 208 -12982
rect 157 -53277 208 -53239
rect 157 -9115 208 -9077
rect 157 -16854 208 -16816
rect 157 -51431 208 -51393
rect 157 -9186 208 -9148
rect 157 -64992 208 -64954
rect 157 -53135 208 -53097
rect 157 -26084 208 -26046
rect 157 -33255 208 -33217
rect 157 -21540 208 -21502
rect 157 -69678 208 -69640
rect 157 -33113 208 -33075
rect 157 -62578 208 -62540
rect 157 -69607 208 -69569
rect 157 -11600 208 -11562
rect 157 -64140 208 -64102
rect 157 -14653 208 -14615
rect 157 -63998 208 -63960
rect 157 -22250 208 -22212
rect 157 -10606 208 -10568
rect 157 -21327 208 -21289
rect 157 -12381 208 -12343
rect 157 -11174 208 -11136
rect 157 -17919 208 -17881
rect 157 -10961 208 -10923
rect 157 -14085 208 -14047
rect 157 -63359 208 -63321
rect 157 -57892 208 -57854
rect 157 -69110 208 -69072
rect 157 -42982 208 -42944
rect 157 -15931 208 -15893
rect 157 -61584 208 -61546
rect 157 -66270 208 -66232
rect 157 -41704 208 -41666
rect 157 -21256 208 -21218
rect 157 -62152 208 -62114
rect 157 -22392 208 -22354
rect 157 -32119 208 -32081
rect 157 -45254 208 -45216
rect 157 -65063 208 -65025
rect 157 -14156 208 -14118
rect 157 -12665 208 -12627
rect 157 -11813 208 -11775
rect 157 -13091 208 -13053
rect 157 -68329 208 -68291
rect 157 -68400 208 -68362
rect 157 -42059 208 -42021
rect 157 -43621 208 -43583
rect 157 -52709 208 -52671
rect 157 -31906 208 -31868
rect 157 -54129 208 -54091
rect 157 -43337 208 -43299
rect 157 -58673 208 -58635
rect 157 -43763 208 -43725
rect 157 -11458 208 -11420
rect 157 -27149 208 -27111
rect 157 -17351 208 -17313
rect 157 -61300 208 -61262
rect 157 -43550 208 -43512
rect 157 -69536 208 -69498
rect 157 -28569 208 -28531
rect 157 -66625 208 -66587
rect 157 -58105 208 -58067
rect 157 -28356 208 -28318
rect 157 -63004 208 -62966
rect 157 -50082 208 -50044
rect 157 -69465 208 -69427
rect 157 -26439 208 -26401
rect 157 -27433 208 -27395
rect 157 -50366 208 -50328
rect 157 -65560 208 -65522
rect 157 -54342 208 -54304
rect 157 -12097 208 -12059
rect 157 -14795 208 -14757
rect 157 -63075 208 -63037
rect 157 -28001 208 -27963
rect 157 -11316 208 -11278
rect 157 -61655 208 -61617
rect 157 -27007 208 -26969
rect 157 -61513 208 -61475
rect 157 -25658 208 -25620
rect 157 -33326 208 -33288
rect 157 -51147 208 -51109
rect 157 -20830 208 -20792
rect 157 -61442 208 -61404
rect 157 -15647 208 -15609
rect 157 -65702 208 -65664
rect 157 -43834 208 -43796
rect 157 -13659 208 -13621
rect 157 -9967 208 -9929
rect 157 -54413 208 -54375
rect 157 -52354 208 -52316
rect 157 -58034 208 -57996
rect 157 -29492 208 -29454
rect 157 -32829 208 -32791
rect 157 -33752 208 -33714
rect 157 -10038 208 -10000
rect 157 -13162 208 -13124
rect 157 -26865 208 -26827
rect 157 -64424 208 -64386
rect 157 -16002 208 -15964
rect 157 -9399 208 -9361
rect 157 -51573 208 -51535
rect 157 -16996 208 -16958
rect 157 -51928 208 -51890
rect 157 -12523 208 -12485
rect 157 -21611 208 -21573
rect 157 -28711 208 -28673
rect 157 -26794 208 -26756
rect 157 -44331 208 -44293
rect 157 -44047 208 -44009
rect 157 -66412 208 -66374
rect 157 -66554 208 -66516
rect 157 -20972 208 -20934
rect 157 -17635 208 -17597
rect 157 -65489 208 -65451
rect 157 -13801 208 -13763
rect 157 -42343 208 -42305
rect 157 -53632 208 -53594
rect 157 -12168 208 -12130
rect 157 -14582 208 -14544
rect 157 -51999 208 -51961
rect 157 -42485 208 -42447
rect 157 -20617 208 -20579
rect 157 -54484 208 -54446
rect 157 -51786 208 -51748
rect 157 -63572 208 -63534
rect 157 -44757 208 -44719
rect 157 -42769 208 -42731
rect 157 -52993 208 -52955
rect -9 -29208 42 -29170
rect -9 -29634 42 -29596
rect -9 -10535 42 -10497
rect -9 -66980 42 -66942
rect -9 -51360 42 -51322
rect -9 -15363 42 -15325
rect -9 -26013 42 -25975
rect -9 -53490 42 -53452
rect -9 -54200 42 -54162
rect -9 -30628 42 -30590
rect -9 -11245 42 -11207
rect -9 -28143 42 -28105
rect -9 -31338 42 -31300
rect -9 -68116 42 -68078
rect -9 -27788 42 -27750
rect -9 -15008 42 -14970
rect -9 -48520 42 -48482
rect -9 -16144 42 -16106
rect -9 -10819 42 -10781
rect -9 -59951 42 -59913
rect -9 -65347 42 -65309
rect -9 -24806 42 -24768
rect -9 -51218 42 -51180
rect -9 -9257 42 -9219
rect -9 -62933 42 -62895
rect -9 -13304 42 -13266
rect -9 -67974 42 -67936
rect -9 -24451 42 -24413
rect -9 -49727 42 -49689
rect -9 -10180 42 -10142
rect -9 -29350 42 -29312
rect -9 -23457 42 -23419
rect -9 -25374 42 -25336
rect -9 -11742 42 -11704
rect -9 -16357 42 -16319
rect -9 -64850 42 -64812
rect -9 -24025 42 -23987
rect -9 -25729 42 -25691
rect -9 -62436 42 -62398
rect -9 -66341 42 -66303
rect -9 -13517 42 -13479
rect -9 -49656 42 -49618
rect -9 -53845 42 -53807
rect -9 -62365 42 -62327
rect -9 -17280 42 -17242
rect -9 -49585 42 -49547
rect -9 -51076 42 -51038
rect -9 -31551 42 -31513
rect -9 -27291 42 -27253
rect -9 -65986 42 -65948
rect -9 -47313 42 -47275
rect -9 -52780 42 -52742
rect -9 -28072 42 -28034
rect -9 -51005 42 -50967
rect -9 -15718 42 -15680
rect -9 -62862 42 -62824
rect -9 -52567 42 -52529
rect -9 -30060 42 -30022
rect -9 -54271 42 -54233
rect -9 -61939 42 -61901
rect -9 -50579 42 -50541
rect -9 -67406 42 -67368
rect -9 -31693 42 -31655
rect -9 -50934 42 -50896
rect -9 -12594 42 -12556
rect -9 -26297 42 -26259
rect -9 -45822 42 -45784
rect -9 -62507 42 -62469
rect -9 -64353 42 -64315
rect -9 -14440 42 -14402
rect -9 -46035 42 -45997
rect -9 -66483 42 -66445
rect -9 -24877 42 -24839
rect -9 -27930 42 -27892
rect -9 -28853 42 -28815
rect -9 -9683 42 -9645
rect -9 -10464 42 -10426
rect -9 -50863 42 -50825
rect -9 -59738 42 -59700
rect -9 -59170 42 -59132
rect -9 -60874 42 -60836
rect -9 -15292 42 -15254
rect -9 -46461 42 -46423
rect -9 -12736 42 -12698
rect -9 -46177 42 -46139
rect -9 -25516 42 -25478
rect -9 -26510 42 -26472
rect -9 -60803 42 -60765
rect -9 -30841 42 -30803
rect -9 -64282 42 -64244
rect -9 -47455 42 -47417
rect -9 -52283 42 -52245
rect -9 -29563 42 -29525
rect -9 -48733 42 -48695
rect -9 -27646 42 -27608
rect -9 -15576 42 -15538
rect -9 -60590 42 -60552
rect -9 -29776 42 -29738
rect -9 -46248 42 -46210
rect -9 -67619 42 -67581
rect -9 -50721 42 -50683
rect -9 -66696 42 -66658
rect -9 -31764 42 -31726
rect -9 -17564 42 -17526
rect -9 -65276 42 -65238
rect -9 -11032 42 -10994
rect -9 -63146 42 -63108
rect -9 -50153 42 -50115
rect -9 -53064 42 -53026
rect -9 -30912 42 -30874
rect -9 -14511 42 -14473
rect -9 -65631 42 -65593
rect -9 -17990 42 -17952
rect -9 -27504 42 -27466
rect -9 -29989 42 -29951
rect -9 -62720 42 -62682
rect -9 -45538 42 -45500
rect -9 -60377 42 -60339
rect -9 -63856 42 -63818
rect -9 -11103 42 -11065
rect -9 -63288 42 -63250
rect -9 -14866 42 -14828
rect -9 -23599 42 -23561
rect -9 -62081 42 -62043
rect -9 -11884 42 -11846
rect -9 -49017 42 -48979
rect -9 -11529 42 -11491
rect -9 -15434 42 -15396
rect -9 -64069 42 -64031
rect -9 -17209 42 -17171
rect -9 -47881 42 -47843
rect -9 -48449 42 -48411
rect -9 -51715 42 -51677
rect -9 -62649 42 -62611
rect -9 -49230 42 -49192
rect -9 -25587 42 -25549
rect -9 -51644 42 -51606
rect -9 -9825 42 -9787
rect -9 -52141 42 -52103
rect -9 -52638 42 -52600
rect -9 -12807 42 -12769
rect -9 -25019 42 -24981
rect -9 -48946 42 -48908
rect -9 -63643 42 -63605
rect -9 -64637 42 -64599
rect -9 -25232 42 -25194
rect -9 -53916 42 -53878
rect -9 -26936 42 -26898
rect -9 -10677 42 -10639
rect -9 -65205 42 -65167
rect -9 -13588 42 -13550
rect -9 -29847 42 -29809
rect -9 -48023 42 -47985
rect -9 -27717 42 -27679
rect -9 -50437 42 -50399
rect -9 -62010 42 -61972
rect -9 -66767 42 -66729
rect -9 -22818 42 -22780
rect -9 -49088 42 -49050
rect -9 -17422 42 -17384
rect -9 -24096 42 -24058
rect -9 -47952 42 -47914
rect -9 -30131 42 -30093
rect -9 -60164 42 -60126
rect -9 -28640 42 -28602
rect -9 -23741 42 -23703
rect -9 -60306 42 -60268
rect -9 -24593 42 -24555
rect -9 -29066 42 -29028
rect -9 -23173 42 -23135
rect -9 -14937 42 -14899
rect -9 -53774 42 -53736
rect -9 -10890 42 -10852
rect -9 -18132 42 -18094
rect -9 -14724 42 -14686
rect -9 -49301 42 -49263
rect -9 -10748 42 -10710
rect -9 -52212 42 -52174
rect -9 -12239 42 -12201
rect -9 -24380 42 -24342
rect -9 -50508 42 -50470
rect -9 -49798 42 -49760
rect -9 -45609 42 -45571
rect -9 -60519 42 -60481
rect -9 -25090 42 -25052
rect -9 -47526 42 -47488
rect -9 -66199 42 -66161
rect -9 -24735 42 -24697
rect -9 -26652 42 -26614
rect -9 -23244 42 -23206
rect -9 -61371 42 -61333
rect -9 -10393 42 -10355
rect -9 -26368 42 -26330
rect -9 -29705 42 -29667
rect -9 -51289 42 -51251
rect -9 -29279 42 -29241
rect -9 -9470 42 -9432
rect -9 -11671 42 -11633
rect -9 -46958 42 -46920
rect -9 -60093 42 -60055
rect -9 -48165 42 -48127
rect -9 -64495 42 -64457
rect -9 -13943 42 -13905
rect -9 -53419 42 -53381
rect -9 -30770 42 -30732
rect -9 -14298 42 -14260
rect -9 -65773 42 -65735
rect -9 -51502 42 -51464
rect -9 -23315 42 -23277
rect -9 -31622 42 -31584
rect -9 -27078 42 -27040
rect -9 -25871 42 -25833
rect -9 -24167 42 -24129
rect -9 -29137 42 -29099
rect -9 -45751 42 -45713
rect -9 -59880 42 -59842
rect -9 -11955 42 -11917
rect -9 -59596 42 -59558
rect -9 -61016 42 -60978
rect -9 -50650 42 -50612
rect -9 -63217 42 -63179
rect -9 -14014 42 -13976
rect -9 -17848 42 -17810
rect -9 -60732 42 -60694
rect -9 -68045 42 -68007
rect -9 -60022 42 -59984
rect -9 -63927 42 -63889
rect -9 -14369 42 -14331
rect -9 -24309 42 -24271
rect -9 -47171 42 -47133
rect -9 -28427 42 -28389
rect -9 -15150 42 -15112
rect -9 -15221 42 -15183
rect -9 -59312 42 -59274
rect -9 -25800 42 -25762
rect -9 -52496 42 -52458
rect -9 -47100 42 -47062
rect -9 -16712 42 -16674
rect -9 -50295 42 -50257
rect -9 -9328 42 -9290
rect -9 -12026 42 -11988
rect -9 -52922 42 -52884
rect -9 -9541 42 -9503
rect -9 -11387 42 -11349
rect -9 -31196 42 -31158
rect -9 -64566 42 -64528
rect -9 -59099 42 -59061
rect -9 -14227 42 -14189
rect -9 -24238 42 -24200
rect -9 -26581 42 -26543
rect -9 -15505 42 -15467
rect -9 -65418 42 -65380
rect -9 -16286 42 -16248
rect -9 -22889 42 -22851
rect -9 -60661 42 -60623
rect -9 -26723 42 -26685
rect -9 -63501 42 -63463
rect -9 -16925 42 -16887
rect -9 -48591 42 -48553
rect -9 -10251 42 -10213
rect -9 -60945 42 -60907
rect -9 -67548 42 -67510
rect -9 -64708 42 -64670
rect -9 -12878 42 -12840
rect -9 -47810 42 -47772
rect -9 -67051 42 -67013
rect -9 -63714 42 -63676
rect -9 -18061 42 -18023
rect -9 -9754 42 -9716
rect -9 -62223 42 -62185
rect -9 -30699 42 -30661
rect -9 -45893 42 -45855
rect -9 -61158 42 -61120
rect -9 -25942 42 -25904
rect -9 -53703 42 -53665
rect -9 -46674 42 -46636
rect -9 -16428 42 -16390
rect -9 -50011 42 -49973
rect -9 -10109 42 -10071
rect -9 -13233 42 -13195
rect -9 -12452 42 -12414
rect -9 -13446 42 -13408
rect -9 -50224 42 -50186
rect -9 -13375 42 -13337
rect -9 -65915 42 -65877
rect -9 -16641 42 -16603
rect -9 -50792 42 -50754
rect -9 -16570 42 -16532
rect -9 -31409 42 -31371
rect -9 -17493 42 -17455
rect -9 -48378 42 -48340
rect -9 -23102 42 -23064
rect -9 -64779 42 -64741
rect -9 -53561 42 -53523
rect -9 -61087 42 -61049
rect -9 -27575 42 -27537
rect -9 -29421 42 -29383
rect -9 -52070 42 -52032
rect -9 -62294 42 -62256
rect -9 -46887 42 -46849
rect -9 -48236 42 -48198
rect -9 -53987 42 -53949
rect -9 -49514 42 -49476
rect -9 -30486 42 -30448
rect -9 -15789 42 -15751
rect -9 -17067 42 -17029
rect -9 -28995 42 -28957
rect -9 -52851 42 -52813
rect -9 -23670 42 -23632
rect -9 -30344 42 -30306
rect -9 -47668 42 -47630
rect -9 -24948 42 -24910
rect -9 -26155 42 -26117
rect -9 -31125 42 -31087
rect -9 -28214 42 -28176
rect -9 -53206 42 -53168
rect -9 -27859 42 -27821
rect -9 -15079 42 -15041
rect -9 -25303 42 -25265
rect -9 -13730 42 -13692
rect -9 -54058 42 -54020
rect -9 -61868 42 -61830
rect -9 -23031 42 -22993
rect -9 -27362 42 -27324
rect -9 -61726 42 -61688
rect -9 -65844 42 -65806
rect -9 -16215 42 -16177
rect -9 -59383 42 -59345
rect -9 -25445 42 -25407
rect -9 -28782 42 -28744
rect -9 -66128 42 -66090
rect -9 -51857 42 -51819
rect -9 -63430 42 -63392
rect -9 -16073 42 -16035
rect -9 -10322 42 -10284
rect -9 -64921 42 -64883
rect -9 -45680 42 -45642
rect -9 -28498 42 -28460
rect -9 -31054 42 -31016
rect -9 -65134 42 -65096
rect -9 -67335 42 -67297
rect -9 -48804 42 -48766
rect -9 -26226 42 -26188
rect -9 -61229 42 -61191
rect -9 -49372 42 -49334
rect -9 -67690 42 -67652
rect -9 -45964 42 -45926
rect -9 -9612 42 -9574
rect -9 -46532 42 -46494
rect -9 -67122 42 -67084
rect -9 -61797 42 -61759
rect -9 -24522 42 -24484
rect -9 -67832 42 -67794
rect -9 -63785 42 -63747
rect -9 -30983 42 -30945
rect -9 -17777 42 -17739
rect -9 -46390 42 -46352
rect -9 -52425 42 -52387
rect -9 -53348 42 -53310
rect -9 -49940 42 -49902
rect -9 -25161 42 -25123
rect -9 -47739 42 -47701
rect -9 -49159 42 -49121
rect -9 -64211 42 -64173
rect -9 -62791 42 -62753
rect -9 -15860 42 -15822
rect -9 -16783 42 -16745
rect -9 -23386 42 -23348
rect -9 -28924 42 -28886
rect -9 -13872 42 -13834
rect -9 -17138 42 -17100
rect -9 -9896 42 -9858
rect -9 -24664 42 -24626
rect -9 -12310 42 -12272
rect -9 -66057 42 -66019
rect -9 -27220 42 -27182
rect -9 -16499 42 -16461
rect -9 -46745 42 -46707
rect -9 -66838 42 -66800
rect -9 -31267 42 -31229
rect -9 -47242 42 -47204
rect -9 -28285 42 -28247
rect -9 -17706 42 -17668
rect -9 -12949 42 -12911
rect -9 -66909 42 -66871
rect -9 -13020 42 -12982
rect -9 -53277 42 -53239
rect -9 -9115 42 -9077
rect -9 -46106 42 -46068
rect -9 -16854 42 -16816
rect -9 -51431 42 -51393
rect -9 -9186 42 -9148
rect -9 -64992 42 -64954
rect -9 -53135 42 -53097
rect -9 -26084 42 -26046
rect -9 -30202 42 -30164
rect -9 -62578 42 -62540
rect -9 -11600 42 -11562
rect -9 -67761 42 -67723
rect -9 -64140 42 -64102
rect -9 -14653 42 -14615
rect -9 -63998 42 -63960
rect -9 -10606 42 -10568
rect -9 -12381 42 -12343
rect -9 -11174 42 -11136
rect -9 -17919 42 -17881
rect -9 -10961 42 -10923
rect -9 -14085 42 -14047
rect -9 -63359 42 -63321
rect -9 -59241 42 -59203
rect -9 -15931 42 -15893
rect -9 -61584 42 -61546
rect -9 -66270 42 -66232
rect -9 -67264 42 -67226
rect -9 -23812 42 -23774
rect -9 -62152 42 -62114
rect -9 -30557 42 -30519
rect -9 -67903 42 -67865
rect -9 -48094 42 -48056
rect -9 -65063 42 -65025
rect -9 -14156 42 -14118
rect -9 -12665 42 -12627
rect -9 -11813 42 -11775
rect -9 -48307 42 -48269
rect -9 -67477 42 -67439
rect -9 -13091 42 -13053
rect -9 -22960 42 -22922
rect -9 -48662 42 -48624
rect -9 -59454 42 -59416
rect -9 -30273 42 -30235
rect -9 -52709 42 -52671
rect -9 -54129 42 -54091
rect -9 -49443 42 -49405
rect -9 -68187 42 -68149
rect -9 -23528 42 -23490
rect -9 -11458 42 -11420
rect -9 -27149 42 -27111
rect -9 -17351 42 -17313
rect -9 -61300 42 -61262
rect -9 -47029 42 -46991
rect -9 -28569 42 -28531
rect -9 -66625 42 -66587
rect -9 -28356 42 -28318
rect -9 -63004 42 -62966
rect -9 -50082 42 -50044
rect -9 -26439 42 -26401
rect -9 -27433 42 -27395
rect -9 -50366 42 -50328
rect -9 -65560 42 -65522
rect -9 -54342 42 -54304
rect -9 -23883 42 -23845
rect -9 -12097 42 -12059
rect -9 -14795 42 -14757
rect -9 -49869 42 -49831
rect -9 -63075 42 -63037
rect -9 -28001 42 -27963
rect -9 -11316 42 -11278
rect -9 -61655 42 -61617
rect -9 -27007 42 -26969
rect -9 -61513 42 -61475
rect -9 -25658 42 -25620
rect -9 -59525 42 -59487
rect -9 -51147 42 -51109
rect -9 -46816 42 -46778
rect -9 -61442 42 -61404
rect -9 -15647 42 -15609
rect -9 -59667 42 -59629
rect -9 -29918 42 -29880
rect -9 -48875 42 -48837
rect -9 -65702 42 -65664
rect -9 -13659 42 -13621
rect -9 -9967 42 -9929
rect -9 -54413 42 -54375
rect -9 -47597 42 -47559
rect -9 -52354 42 -52316
rect -9 -29492 42 -29454
rect -9 -10038 42 -10000
rect -9 -30415 42 -30377
rect -9 -60235 42 -60197
rect -9 -13162 42 -13124
rect -9 -26865 42 -26827
rect -9 -64424 42 -64386
rect -9 -16002 42 -15964
rect -9 -47384 42 -47346
rect -9 -9399 42 -9361
rect -9 -51573 42 -51535
rect -9 -16996 42 -16958
rect -9 -51928 42 -51890
rect -9 -12523 42 -12485
rect -9 -31480 42 -31442
rect -9 -28711 42 -28673
rect -9 -26794 42 -26756
rect -9 -66412 42 -66374
rect -9 -23954 42 -23916
rect -9 -66554 42 -66516
rect -9 -17635 42 -17597
rect -9 -59809 42 -59771
rect -9 -65489 42 -65451
rect -9 -13801 42 -13763
rect -9 -60448 42 -60410
rect -9 -53632 42 -53594
rect -9 -12168 42 -12130
rect -9 -14582 42 -14544
rect -9 -46319 42 -46281
rect -9 -51999 42 -51961
rect -9 -67193 42 -67155
rect -9 -54484 42 -54446
rect -9 -51786 42 -51748
rect -9 -63572 42 -63534
rect -9 -46603 42 -46565
rect -9 -52993 42 -52955
<< pdiff >>
rect 904 138 955 227
rect 738 138 789 227
rect 655 138 706 227
rect 489 138 540 227
rect 406 138 457 227
rect 240 138 291 227
rect 157 138 208 227
rect -9 138 42 227
<< ndiffc >>
<< pdiffc >>
rect 921 146 938 163
rect 912 202 947 219
rect 755 146 772 163
rect 746 202 781 219
rect 672 146 689 163
rect 663 202 698 219
rect 506 146 523 163
rect 497 202 532 219
rect 423 146 440 163
rect 414 202 449 219
rect 257 146 274 163
rect 248 202 283 219
rect 174 146 191 163
rect 165 202 200 219
rect 8 146 25 163
rect -1 202 34 219
<< psubdiff >>
rect -27 79 973 107
<< nsubdiff >>
rect -9 254 955 282
<< psubdiffcont >>
rect -15 79 961 107
<< nsubdiffcont >>
rect 3 254 943 282
<< ndcontact >>
rect 838 -9140 855 -9123
rect 340 -9140 357 -9123
rect 91 -9140 108 -9123
rect 589 -9140 606 -9123
rect 838 -9282 855 -9265
rect 340 -9282 357 -9265
rect 91 -9282 108 -9265
rect 589 -9282 606 -9265
rect 838 -9424 855 -9407
rect 340 -9424 357 -9407
rect 91 -9424 108 -9407
rect 589 -9424 606 -9407
rect 838 -9566 855 -9549
rect 340 -9566 357 -9549
rect 91 -9566 108 -9549
rect 589 -9566 606 -9549
rect 838 -9708 855 -9691
rect 340 -9708 357 -9691
rect 91 -9708 108 -9691
rect 589 -9708 606 -9691
rect 838 -9850 855 -9833
rect 340 -9850 357 -9833
rect 91 -9850 108 -9833
rect 589 -9850 606 -9833
rect 838 -9992 855 -9975
rect 340 -9992 357 -9975
rect 91 -9992 108 -9975
rect 589 -9992 606 -9975
rect 838 -10134 855 -10117
rect 340 -10134 357 -10117
rect 91 -10134 108 -10117
rect 589 -10134 606 -10117
rect 838 -10276 855 -10259
rect 340 -10276 357 -10259
rect 91 -10276 108 -10259
rect 589 -10276 606 -10259
rect 838 -10418 855 -10401
rect 340 -10418 357 -10401
rect 91 -10418 108 -10401
rect 589 -10418 606 -10401
rect 838 -10560 855 -10543
rect 340 -10560 357 -10543
rect 91 -10560 108 -10543
rect 589 -10560 606 -10543
rect 838 -10702 855 -10685
rect 340 -10702 357 -10685
rect 91 -10702 108 -10685
rect 589 -10702 606 -10685
rect 838 -10844 855 -10827
rect 340 -10844 357 -10827
rect 91 -10844 108 -10827
rect 589 -10844 606 -10827
rect 838 -10986 855 -10969
rect 340 -10986 357 -10969
rect 91 -10986 108 -10969
rect 589 -10986 606 -10969
rect 838 -11128 855 -11111
rect 340 -11128 357 -11111
rect 91 -11128 108 -11111
rect 589 -11128 606 -11111
rect 838 -11270 855 -11253
rect 340 -11270 357 -11253
rect 91 -11270 108 -11253
rect 589 -11270 606 -11253
rect 838 -11412 855 -11395
rect 340 -11412 357 -11395
rect 91 -11412 108 -11395
rect 589 -11412 606 -11395
rect 838 -11554 855 -11537
rect 340 -11554 357 -11537
rect 91 -11554 108 -11537
rect 589 -11554 606 -11537
rect 838 -11696 855 -11679
rect 340 -11696 357 -11679
rect 91 -11696 108 -11679
rect 589 -11696 606 -11679
rect 838 -11838 855 -11821
rect 340 -11838 357 -11821
rect 91 -11838 108 -11821
rect 589 -11838 606 -11821
rect 838 -11980 855 -11963
rect 340 -11980 357 -11963
rect 91 -11980 108 -11963
rect 589 -11980 606 -11963
rect 838 -12122 855 -12105
rect 340 -12122 357 -12105
rect 91 -12122 108 -12105
rect 589 -12122 606 -12105
rect 838 -12264 855 -12247
rect 340 -12264 357 -12247
rect 91 -12264 108 -12247
rect 589 -12264 606 -12247
rect 838 -12406 855 -12389
rect 340 -12406 357 -12389
rect 91 -12406 108 -12389
rect 589 -12406 606 -12389
rect 838 -12548 855 -12531
rect 340 -12548 357 -12531
rect 91 -12548 108 -12531
rect 589 -12548 606 -12531
rect 838 -12690 855 -12673
rect 340 -12690 357 -12673
rect 91 -12690 108 -12673
rect 589 -12690 606 -12673
rect 838 -12832 855 -12815
rect 340 -12832 357 -12815
rect 91 -12832 108 -12815
rect 589 -12832 606 -12815
rect 838 -12974 855 -12957
rect 340 -12974 357 -12957
rect 91 -12974 108 -12957
rect 589 -12974 606 -12957
rect 838 -13116 855 -13099
rect 340 -13116 357 -13099
rect 91 -13116 108 -13099
rect 589 -13116 606 -13099
rect 838 -13258 855 -13241
rect 340 -13258 357 -13241
rect 91 -13258 108 -13241
rect 589 -13258 606 -13241
rect 838 -13400 855 -13383
rect 340 -13400 357 -13383
rect 91 -13400 108 -13383
rect 589 -13400 606 -13383
rect 838 -13542 855 -13525
rect 340 -13542 357 -13525
rect 91 -13542 108 -13525
rect 589 -13542 606 -13525
rect 838 -13684 855 -13667
rect 340 -13684 357 -13667
rect 91 -13684 108 -13667
rect 589 -13684 606 -13667
rect 838 -13826 855 -13809
rect 340 -13826 357 -13809
rect 91 -13826 108 -13809
rect 589 -13826 606 -13809
rect 838 -13968 855 -13951
rect 340 -13968 357 -13951
rect 91 -13968 108 -13951
rect 589 -13968 606 -13951
rect 838 -14110 855 -14093
rect 340 -14110 357 -14093
rect 91 -14110 108 -14093
rect 589 -14110 606 -14093
rect 838 -14252 855 -14235
rect 340 -14252 357 -14235
rect 91 -14252 108 -14235
rect 589 -14252 606 -14235
rect 838 -14394 855 -14377
rect 340 -14394 357 -14377
rect 91 -14394 108 -14377
rect 589 -14394 606 -14377
rect 838 -14536 855 -14519
rect 340 -14536 357 -14519
rect 91 -14536 108 -14519
rect 589 -14536 606 -14519
rect 838 -14678 855 -14661
rect 340 -14678 357 -14661
rect 91 -14678 108 -14661
rect 589 -14678 606 -14661
rect 838 -14820 855 -14803
rect 340 -14820 357 -14803
rect 91 -14820 108 -14803
rect 589 -14820 606 -14803
rect 838 -14962 855 -14945
rect 340 -14962 357 -14945
rect 91 -14962 108 -14945
rect 589 -14962 606 -14945
rect 838 -15104 855 -15087
rect 340 -15104 357 -15087
rect 91 -15104 108 -15087
rect 589 -15104 606 -15087
rect 838 -15246 855 -15229
rect 340 -15246 357 -15229
rect 91 -15246 108 -15229
rect 589 -15246 606 -15229
rect 838 -15388 855 -15371
rect 340 -15388 357 -15371
rect 91 -15388 108 -15371
rect 589 -15388 606 -15371
rect 838 -15530 855 -15513
rect 340 -15530 357 -15513
rect 91 -15530 108 -15513
rect 589 -15530 606 -15513
rect 838 -15672 855 -15655
rect 340 -15672 357 -15655
rect 91 -15672 108 -15655
rect 589 -15672 606 -15655
rect 838 -15814 855 -15797
rect 340 -15814 357 -15797
rect 91 -15814 108 -15797
rect 589 -15814 606 -15797
rect 838 -15956 855 -15939
rect 340 -15956 357 -15939
rect 91 -15956 108 -15939
rect 589 -15956 606 -15939
rect 838 -16098 855 -16081
rect 340 -16098 357 -16081
rect 91 -16098 108 -16081
rect 589 -16098 606 -16081
rect 838 -16240 855 -16223
rect 340 -16240 357 -16223
rect 91 -16240 108 -16223
rect 589 -16240 606 -16223
rect 838 -16382 855 -16365
rect 340 -16382 357 -16365
rect 91 -16382 108 -16365
rect 589 -16382 606 -16365
rect 838 -16524 855 -16507
rect 340 -16524 357 -16507
rect 91 -16524 108 -16507
rect 589 -16524 606 -16507
rect 838 -16666 855 -16649
rect 340 -16666 357 -16649
rect 91 -16666 108 -16649
rect 589 -16666 606 -16649
rect 838 -16808 855 -16791
rect 340 -16808 357 -16791
rect 91 -16808 108 -16791
rect 589 -16808 606 -16791
rect 838 -16950 855 -16933
rect 340 -16950 357 -16933
rect 91 -16950 108 -16933
rect 589 -16950 606 -16933
rect 838 -17092 855 -17075
rect 340 -17092 357 -17075
rect 91 -17092 108 -17075
rect 589 -17092 606 -17075
rect 838 -17234 855 -17217
rect 340 -17234 357 -17217
rect 91 -17234 108 -17217
rect 589 -17234 606 -17217
rect 838 -17376 855 -17359
rect 340 -17376 357 -17359
rect 91 -17376 108 -17359
rect 589 -17376 606 -17359
rect 838 -17518 855 -17501
rect 340 -17518 357 -17501
rect 91 -17518 108 -17501
rect 589 -17518 606 -17501
rect 838 -17660 855 -17643
rect 340 -17660 357 -17643
rect 91 -17660 108 -17643
rect 589 -17660 606 -17643
rect 838 -17802 855 -17785
rect 340 -17802 357 -17785
rect 91 -17802 108 -17785
rect 589 -17802 606 -17785
rect 838 -17944 855 -17927
rect 340 -17944 357 -17927
rect 91 -17944 108 -17927
rect 589 -17944 606 -17927
rect 838 -18086 855 -18069
rect 340 -18086 357 -18069
rect 91 -18086 108 -18069
rect 589 -18086 606 -18069
rect 838 -18228 855 -18211
rect 838 -18370 855 -18353
rect 589 -18370 606 -18353
rect 838 -18512 855 -18495
rect 589 -18512 606 -18495
rect 838 -18654 855 -18637
rect 589 -18654 606 -18637
rect 838 -18796 855 -18779
rect 340 -18796 357 -18779
rect 589 -18796 606 -18779
rect 838 -18938 855 -18921
rect 340 -18938 357 -18921
rect 589 -18938 606 -18921
rect 838 -19080 855 -19063
rect 340 -19080 357 -19063
rect 589 -19080 606 -19063
rect 838 -19222 855 -19205
rect 340 -19222 357 -19205
rect 589 -19222 606 -19205
rect 838 -19364 855 -19347
rect 340 -19364 357 -19347
rect 589 -19364 606 -19347
rect 838 -19506 855 -19489
rect 340 -19506 357 -19489
rect 589 -19506 606 -19489
rect 838 -19648 855 -19631
rect 340 -19648 357 -19631
rect 589 -19648 606 -19631
rect 838 -19790 855 -19773
rect 340 -19790 357 -19773
rect 589 -19790 606 -19773
rect 838 -19932 855 -19915
rect 340 -19932 357 -19915
rect 589 -19932 606 -19915
rect 838 -20074 855 -20057
rect 340 -20074 357 -20057
rect 589 -20074 606 -20057
rect 838 -20216 855 -20199
rect 340 -20216 357 -20199
rect 589 -20216 606 -20199
rect 838 -20358 855 -20341
rect 340 -20358 357 -20341
rect 589 -20358 606 -20341
rect 838 -20500 855 -20483
rect 340 -20500 357 -20483
rect 91 -20500 108 -20483
rect 589 -20500 606 -20483
rect 838 -20642 855 -20625
rect 91 -20642 108 -20625
rect 589 -20642 606 -20625
rect 838 -20784 855 -20767
rect 91 -20784 108 -20767
rect 589 -20784 606 -20767
rect 838 -20926 855 -20909
rect 91 -20926 108 -20909
rect 589 -20926 606 -20909
rect 838 -21068 855 -21051
rect 340 -21068 357 -21051
rect 91 -21068 108 -21051
rect 589 -21068 606 -21051
rect 838 -21210 855 -21193
rect 340 -21210 357 -21193
rect 91 -21210 108 -21193
rect 589 -21210 606 -21193
rect 838 -21352 855 -21335
rect 340 -21352 357 -21335
rect 91 -21352 108 -21335
rect 589 -21352 606 -21335
rect 838 -21494 855 -21477
rect 340 -21494 357 -21477
rect 91 -21494 108 -21477
rect 589 -21494 606 -21477
rect 838 -21636 855 -21619
rect 340 -21636 357 -21619
rect 91 -21636 108 -21619
rect 589 -21636 606 -21619
rect 838 -21778 855 -21761
rect 340 -21778 357 -21761
rect 91 -21778 108 -21761
rect 589 -21778 606 -21761
rect 838 -21920 855 -21903
rect 340 -21920 357 -21903
rect 91 -21920 108 -21903
rect 589 -21920 606 -21903
rect 838 -22062 855 -22045
rect 340 -22062 357 -22045
rect 91 -22062 108 -22045
rect 589 -22062 606 -22045
rect 838 -22204 855 -22187
rect 340 -22204 357 -22187
rect 91 -22204 108 -22187
rect 589 -22204 606 -22187
rect 838 -22346 855 -22329
rect 340 -22346 357 -22329
rect 91 -22346 108 -22329
rect 589 -22346 606 -22329
rect 838 -22488 855 -22471
rect 340 -22488 357 -22471
rect 91 -22488 108 -22471
rect 589 -22488 606 -22471
rect 838 -22630 855 -22613
rect 340 -22630 357 -22613
rect 91 -22630 108 -22613
rect 589 -22630 606 -22613
rect 838 -22772 855 -22755
rect 340 -22772 357 -22755
rect 91 -22772 108 -22755
rect 589 -22772 606 -22755
rect 838 -22914 855 -22897
rect 91 -22914 108 -22897
rect 589 -22914 606 -22897
rect 838 -23056 855 -23039
rect 91 -23056 108 -23039
rect 589 -23056 606 -23039
rect 838 -23198 855 -23181
rect 91 -23198 108 -23181
rect 589 -23198 606 -23181
rect 838 -23340 855 -23323
rect 340 -23340 357 -23323
rect 91 -23340 108 -23323
rect 589 -23340 606 -23323
rect 838 -23482 855 -23465
rect 340 -23482 357 -23465
rect 91 -23482 108 -23465
rect 589 -23482 606 -23465
rect 838 -23624 855 -23607
rect 340 -23624 357 -23607
rect 91 -23624 108 -23607
rect 589 -23624 606 -23607
rect 838 -23766 855 -23749
rect 340 -23766 357 -23749
rect 91 -23766 108 -23749
rect 589 -23766 606 -23749
rect 838 -23908 855 -23891
rect 340 -23908 357 -23891
rect 91 -23908 108 -23891
rect 589 -23908 606 -23891
rect 838 -24050 855 -24033
rect 340 -24050 357 -24033
rect 91 -24050 108 -24033
rect 589 -24050 606 -24033
rect 838 -24192 855 -24175
rect 340 -24192 357 -24175
rect 91 -24192 108 -24175
rect 589 -24192 606 -24175
rect 838 -24334 855 -24317
rect 340 -24334 357 -24317
rect 91 -24334 108 -24317
rect 589 -24334 606 -24317
rect 838 -24476 855 -24459
rect 340 -24476 357 -24459
rect 91 -24476 108 -24459
rect 589 -24476 606 -24459
rect 838 -24618 855 -24601
rect 340 -24618 357 -24601
rect 91 -24618 108 -24601
rect 589 -24618 606 -24601
rect 838 -24760 855 -24743
rect 340 -24760 357 -24743
rect 91 -24760 108 -24743
rect 589 -24760 606 -24743
rect 838 -24902 855 -24885
rect 340 -24902 357 -24885
rect 91 -24902 108 -24885
rect 589 -24902 606 -24885
rect 838 -25044 855 -25027
rect 340 -25044 357 -25027
rect 91 -25044 108 -25027
rect 589 -25044 606 -25027
rect 838 -25186 855 -25169
rect 91 -25186 108 -25169
rect 589 -25186 606 -25169
rect 838 -25328 855 -25311
rect 91 -25328 108 -25311
rect 589 -25328 606 -25311
rect 838 -25470 855 -25453
rect 91 -25470 108 -25453
rect 589 -25470 606 -25453
rect 838 -25612 855 -25595
rect 340 -25612 357 -25595
rect 91 -25612 108 -25595
rect 589 -25612 606 -25595
rect 838 -25754 855 -25737
rect 340 -25754 357 -25737
rect 91 -25754 108 -25737
rect 589 -25754 606 -25737
rect 838 -25896 855 -25879
rect 340 -25896 357 -25879
rect 91 -25896 108 -25879
rect 589 -25896 606 -25879
rect 838 -26038 855 -26021
rect 340 -26038 357 -26021
rect 91 -26038 108 -26021
rect 589 -26038 606 -26021
rect 838 -26180 855 -26163
rect 340 -26180 357 -26163
rect 91 -26180 108 -26163
rect 589 -26180 606 -26163
rect 838 -26322 855 -26305
rect 340 -26322 357 -26305
rect 91 -26322 108 -26305
rect 589 -26322 606 -26305
rect 838 -26464 855 -26447
rect 340 -26464 357 -26447
rect 91 -26464 108 -26447
rect 589 -26464 606 -26447
rect 838 -26606 855 -26589
rect 340 -26606 357 -26589
rect 91 -26606 108 -26589
rect 589 -26606 606 -26589
rect 838 -26748 855 -26731
rect 340 -26748 357 -26731
rect 91 -26748 108 -26731
rect 589 -26748 606 -26731
rect 838 -26890 855 -26873
rect 340 -26890 357 -26873
rect 91 -26890 108 -26873
rect 589 -26890 606 -26873
rect 838 -27032 855 -27015
rect 340 -27032 357 -27015
rect 91 -27032 108 -27015
rect 589 -27032 606 -27015
rect 838 -27174 855 -27157
rect 340 -27174 357 -27157
rect 91 -27174 108 -27157
rect 589 -27174 606 -27157
rect 838 -27316 855 -27299
rect 340 -27316 357 -27299
rect 91 -27316 108 -27299
rect 589 -27316 606 -27299
rect 838 -27458 855 -27441
rect 340 -27458 357 -27441
rect 91 -27458 108 -27441
rect 589 -27458 606 -27441
rect 838 -27600 855 -27583
rect 340 -27600 357 -27583
rect 91 -27600 108 -27583
rect 589 -27600 606 -27583
rect 838 -27742 855 -27725
rect 340 -27742 357 -27725
rect 91 -27742 108 -27725
rect 838 -27884 855 -27867
rect 340 -27884 357 -27867
rect 91 -27884 108 -27867
rect 589 -27884 606 -27867
rect 838 -28026 855 -28009
rect 340 -28026 357 -28009
rect 91 -28026 108 -28009
rect 589 -28026 606 -28009
rect 838 -28168 855 -28151
rect 340 -28168 357 -28151
rect 91 -28168 108 -28151
rect 589 -28168 606 -28151
rect 838 -28310 855 -28293
rect 340 -28310 357 -28293
rect 91 -28310 108 -28293
rect 838 -28452 855 -28435
rect 340 -28452 357 -28435
rect 91 -28452 108 -28435
rect 589 -28452 606 -28435
rect 838 -28594 855 -28577
rect 340 -28594 357 -28577
rect 91 -28594 108 -28577
rect 589 -28594 606 -28577
rect 838 -28736 855 -28719
rect 340 -28736 357 -28719
rect 91 -28736 108 -28719
rect 589 -28736 606 -28719
rect 838 -28878 855 -28861
rect 340 -28878 357 -28861
rect 91 -28878 108 -28861
rect 838 -29020 855 -29003
rect 91 -29020 108 -29003
rect 589 -29020 606 -29003
rect 838 -29162 855 -29145
rect 91 -29162 108 -29145
rect 589 -29162 606 -29145
rect 838 -29304 855 -29287
rect 91 -29304 108 -29287
rect 589 -29304 606 -29287
rect 838 -29446 855 -29429
rect 91 -29446 108 -29429
rect 838 -29588 855 -29571
rect 340 -29588 357 -29571
rect 91 -29588 108 -29571
rect 589 -29588 606 -29571
rect 838 -29730 855 -29713
rect 340 -29730 357 -29713
rect 91 -29730 108 -29713
rect 589 -29730 606 -29713
rect 838 -29872 855 -29855
rect 340 -29872 357 -29855
rect 91 -29872 108 -29855
rect 589 -29872 606 -29855
rect 838 -30014 855 -29997
rect 340 -30014 357 -29997
rect 91 -30014 108 -29997
rect 838 -30156 855 -30139
rect 340 -30156 357 -30139
rect 91 -30156 108 -30139
rect 589 -30156 606 -30139
rect 838 -30298 855 -30281
rect 340 -30298 357 -30281
rect 91 -30298 108 -30281
rect 589 -30298 606 -30281
rect 838 -30440 855 -30423
rect 340 -30440 357 -30423
rect 91 -30440 108 -30423
rect 589 -30440 606 -30423
rect 838 -30582 855 -30565
rect 340 -30582 357 -30565
rect 91 -30582 108 -30565
rect 838 -30724 855 -30707
rect 340 -30724 357 -30707
rect 91 -30724 108 -30707
rect 589 -30724 606 -30707
rect 838 -30866 855 -30849
rect 340 -30866 357 -30849
rect 91 -30866 108 -30849
rect 589 -30866 606 -30849
rect 838 -31008 855 -30991
rect 340 -31008 357 -30991
rect 91 -31008 108 -30991
rect 589 -31008 606 -30991
rect 838 -31150 855 -31133
rect 340 -31150 357 -31133
rect 91 -31150 108 -31133
rect 838 -31292 855 -31275
rect 91 -31292 108 -31275
rect 589 -31292 606 -31275
rect 838 -31434 855 -31417
rect 91 -31434 108 -31417
rect 589 -31434 606 -31417
rect 838 -31576 855 -31559
rect 91 -31576 108 -31559
rect 589 -31576 606 -31559
rect 838 -31718 855 -31701
rect 91 -31718 108 -31701
rect 838 -31860 855 -31843
rect 340 -31860 357 -31843
rect 91 -31860 108 -31843
rect 589 -31860 606 -31843
rect 838 -32002 855 -31985
rect 340 -32002 357 -31985
rect 91 -32002 108 -31985
rect 589 -32002 606 -31985
rect 838 -32144 855 -32127
rect 340 -32144 357 -32127
rect 91 -32144 108 -32127
rect 589 -32144 606 -32127
rect 838 -32286 855 -32269
rect 340 -32286 357 -32269
rect 91 -32286 108 -32269
rect 838 -32428 855 -32411
rect 340 -32428 357 -32411
rect 91 -32428 108 -32411
rect 589 -32428 606 -32411
rect 838 -32570 855 -32553
rect 340 -32570 357 -32553
rect 91 -32570 108 -32553
rect 589 -32570 606 -32553
rect 838 -32712 855 -32695
rect 340 -32712 357 -32695
rect 91 -32712 108 -32695
rect 589 -32712 606 -32695
rect 838 -32854 855 -32837
rect 340 -32854 357 -32837
rect 91 -32854 108 -32837
rect 838 -32996 855 -32979
rect 340 -32996 357 -32979
rect 91 -32996 108 -32979
rect 589 -32996 606 -32979
rect 838 -33138 855 -33121
rect 340 -33138 357 -33121
rect 91 -33138 108 -33121
rect 589 -33138 606 -33121
rect 838 -33280 855 -33263
rect 340 -33280 357 -33263
rect 91 -33280 108 -33263
rect 589 -33280 606 -33263
rect 838 -33422 855 -33405
rect 340 -33422 357 -33405
rect 91 -33422 108 -33405
rect 838 -33564 855 -33547
rect 91 -33564 108 -33547
rect 589 -33564 606 -33547
rect 838 -33706 855 -33689
rect 91 -33706 108 -33689
rect 589 -33706 606 -33689
rect 838 -33848 855 -33831
rect 91 -33848 108 -33831
rect 589 -33848 606 -33831
rect 838 -33990 855 -33973
rect 91 -33990 108 -33973
rect 838 -34132 855 -34115
rect 340 -34132 357 -34115
rect 589 -34132 606 -34115
rect 838 -34274 855 -34257
rect 340 -34274 357 -34257
rect 589 -34274 606 -34257
rect 838 -34416 855 -34399
rect 340 -34416 357 -34399
rect 589 -34416 606 -34399
rect 838 -34558 855 -34541
rect 340 -34558 357 -34541
rect 838 -34700 855 -34683
rect 340 -34700 357 -34683
rect 589 -34700 606 -34683
rect 838 -34842 855 -34825
rect 340 -34842 357 -34825
rect 589 -34842 606 -34825
rect 838 -34984 855 -34967
rect 340 -34984 357 -34967
rect 589 -34984 606 -34967
rect 838 -35126 855 -35109
rect 340 -35126 357 -35109
rect 838 -35268 855 -35251
rect 340 -35268 357 -35251
rect 589 -35268 606 -35251
rect 838 -35410 855 -35393
rect 340 -35410 357 -35393
rect 589 -35410 606 -35393
rect 838 -35552 855 -35535
rect 340 -35552 357 -35535
rect 589 -35552 606 -35535
rect 838 -35694 855 -35677
rect 340 -35694 357 -35677
rect 838 -35836 855 -35819
rect 589 -35836 606 -35819
rect 838 -35978 855 -35961
rect 589 -35978 606 -35961
rect 838 -36120 855 -36103
rect 589 -36120 606 -36103
rect 838 -36262 855 -36245
rect 838 -36546 855 -36529
rect 838 -36688 855 -36671
rect 589 -36688 606 -36671
rect 838 -36830 855 -36813
rect 589 -36830 606 -36813
rect 838 -36972 855 -36955
rect 589 -36972 606 -36955
rect 838 -37114 855 -37097
rect 589 -37114 606 -37097
rect 838 -37256 855 -37239
rect 589 -37256 606 -37239
rect 838 -37398 855 -37381
rect 589 -37398 606 -37381
rect 838 -37540 855 -37523
rect 340 -37540 357 -37523
rect 589 -37540 606 -37523
rect 838 -37682 855 -37665
rect 340 -37682 357 -37665
rect 838 -37824 855 -37807
rect 340 -37824 357 -37807
rect 589 -37824 606 -37807
rect 838 -37966 855 -37949
rect 340 -37966 357 -37949
rect 589 -37966 606 -37949
rect 838 -38108 855 -38091
rect 340 -38108 357 -38091
rect 589 -38108 606 -38091
rect 838 -38250 855 -38233
rect 340 -38250 357 -38233
rect 589 -38250 606 -38233
rect 838 -38392 855 -38375
rect 340 -38392 357 -38375
rect 589 -38392 606 -38375
rect 838 -38534 855 -38517
rect 340 -38534 357 -38517
rect 589 -38534 606 -38517
rect 838 -38676 855 -38659
rect 340 -38676 357 -38659
rect 589 -38676 606 -38659
rect 838 -38818 855 -38801
rect 340 -38818 357 -38801
rect 838 -38960 855 -38943
rect 340 -38960 357 -38943
rect 589 -38960 606 -38943
rect 838 -39102 855 -39085
rect 340 -39102 357 -39085
rect 589 -39102 606 -39085
rect 838 -39244 855 -39227
rect 340 -39244 357 -39227
rect 589 -39244 606 -39227
rect 838 -39386 855 -39369
rect 340 -39386 357 -39369
rect 589 -39386 606 -39369
rect 838 -39528 855 -39511
rect 340 -39528 357 -39511
rect 589 -39528 606 -39511
rect 838 -39670 855 -39653
rect 340 -39670 357 -39653
rect 589 -39670 606 -39653
rect 838 -39812 855 -39795
rect 340 -39812 357 -39795
rect 589 -39812 606 -39795
rect 838 -39954 855 -39937
rect 340 -39954 357 -39937
rect 838 -40096 855 -40079
rect 340 -40096 357 -40079
rect 589 -40096 606 -40079
rect 838 -40238 855 -40221
rect 340 -40238 357 -40221
rect 589 -40238 606 -40221
rect 838 -40380 855 -40363
rect 340 -40380 357 -40363
rect 589 -40380 606 -40363
rect 838 -40522 855 -40505
rect 340 -40522 357 -40505
rect 589 -40522 606 -40505
rect 838 -40664 855 -40647
rect 340 -40664 357 -40647
rect 589 -40664 606 -40647
rect 838 -40806 855 -40789
rect 340 -40806 357 -40789
rect 589 -40806 606 -40789
rect 838 -40948 855 -40931
rect 340 -40948 357 -40931
rect 91 -40948 108 -40931
rect 589 -40948 606 -40931
rect 838 -41090 855 -41073
rect 91 -41090 108 -41073
rect 838 -41232 855 -41215
rect 91 -41232 108 -41215
rect 589 -41232 606 -41215
rect 838 -41374 855 -41357
rect 91 -41374 108 -41357
rect 589 -41374 606 -41357
rect 838 -41516 855 -41499
rect 91 -41516 108 -41499
rect 589 -41516 606 -41499
rect 838 -41658 855 -41641
rect 91 -41658 108 -41641
rect 589 -41658 606 -41641
rect 838 -41800 855 -41783
rect 91 -41800 108 -41783
rect 589 -41800 606 -41783
rect 838 -41942 855 -41925
rect 91 -41942 108 -41925
rect 589 -41942 606 -41925
rect 838 -42084 855 -42067
rect 340 -42084 357 -42067
rect 91 -42084 108 -42067
rect 589 -42084 606 -42067
rect 838 -42226 855 -42209
rect 340 -42226 357 -42209
rect 91 -42226 108 -42209
rect 838 -42368 855 -42351
rect 340 -42368 357 -42351
rect 91 -42368 108 -42351
rect 589 -42368 606 -42351
rect 838 -42510 855 -42493
rect 340 -42510 357 -42493
rect 91 -42510 108 -42493
rect 589 -42510 606 -42493
rect 838 -42652 855 -42635
rect 340 -42652 357 -42635
rect 91 -42652 108 -42635
rect 589 -42652 606 -42635
rect 838 -42794 855 -42777
rect 340 -42794 357 -42777
rect 91 -42794 108 -42777
rect 589 -42794 606 -42777
rect 838 -42936 855 -42919
rect 340 -42936 357 -42919
rect 91 -42936 108 -42919
rect 589 -42936 606 -42919
rect 838 -43078 855 -43061
rect 340 -43078 357 -43061
rect 91 -43078 108 -43061
rect 589 -43078 606 -43061
rect 838 -43220 855 -43203
rect 340 -43220 357 -43203
rect 91 -43220 108 -43203
rect 589 -43220 606 -43203
rect 838 -43362 855 -43345
rect 340 -43362 357 -43345
rect 91 -43362 108 -43345
rect 838 -43504 855 -43487
rect 340 -43504 357 -43487
rect 91 -43504 108 -43487
rect 589 -43504 606 -43487
rect 838 -43646 855 -43629
rect 340 -43646 357 -43629
rect 91 -43646 108 -43629
rect 589 -43646 606 -43629
rect 838 -43788 855 -43771
rect 340 -43788 357 -43771
rect 91 -43788 108 -43771
rect 589 -43788 606 -43771
rect 838 -43930 855 -43913
rect 340 -43930 357 -43913
rect 91 -43930 108 -43913
rect 589 -43930 606 -43913
rect 838 -44072 855 -44055
rect 340 -44072 357 -44055
rect 91 -44072 108 -44055
rect 589 -44072 606 -44055
rect 838 -44214 855 -44197
rect 340 -44214 357 -44197
rect 91 -44214 108 -44197
rect 589 -44214 606 -44197
rect 838 -44356 855 -44339
rect 340 -44356 357 -44339
rect 91 -44356 108 -44339
rect 589 -44356 606 -44339
rect 838 -44498 855 -44481
rect 340 -44498 357 -44481
rect 91 -44498 108 -44481
rect 838 -44640 855 -44623
rect 340 -44640 357 -44623
rect 91 -44640 108 -44623
rect 589 -44640 606 -44623
rect 838 -44782 855 -44765
rect 340 -44782 357 -44765
rect 91 -44782 108 -44765
rect 589 -44782 606 -44765
rect 838 -44924 855 -44907
rect 340 -44924 357 -44907
rect 91 -44924 108 -44907
rect 589 -44924 606 -44907
rect 838 -45066 855 -45049
rect 340 -45066 357 -45049
rect 91 -45066 108 -45049
rect 589 -45066 606 -45049
rect 838 -45208 855 -45191
rect 340 -45208 357 -45191
rect 91 -45208 108 -45191
rect 589 -45208 606 -45191
rect 838 -45350 855 -45333
rect 340 -45350 357 -45333
rect 91 -45350 108 -45333
rect 589 -45350 606 -45333
rect 838 -45492 855 -45475
rect 340 -45492 357 -45475
rect 91 -45492 108 -45475
rect 589 -45492 606 -45475
rect 838 -45634 855 -45617
rect 91 -45634 108 -45617
rect 838 -45776 855 -45759
rect 91 -45776 108 -45759
rect 589 -45776 606 -45759
rect 838 -45918 855 -45901
rect 91 -45918 108 -45901
rect 589 -45918 606 -45901
rect 838 -46060 855 -46043
rect 91 -46060 108 -46043
rect 589 -46060 606 -46043
rect 838 -46202 855 -46185
rect 91 -46202 108 -46185
rect 589 -46202 606 -46185
rect 838 -46344 855 -46327
rect 91 -46344 108 -46327
rect 589 -46344 606 -46327
rect 838 -46486 855 -46469
rect 91 -46486 108 -46469
rect 589 -46486 606 -46469
rect 838 -46628 855 -46611
rect 340 -46628 357 -46611
rect 91 -46628 108 -46611
rect 589 -46628 606 -46611
rect 838 -46770 855 -46753
rect 340 -46770 357 -46753
rect 91 -46770 108 -46753
rect 838 -46912 855 -46895
rect 340 -46912 357 -46895
rect 91 -46912 108 -46895
rect 589 -46912 606 -46895
rect 838 -47054 855 -47037
rect 340 -47054 357 -47037
rect 91 -47054 108 -47037
rect 589 -47054 606 -47037
rect 838 -47196 855 -47179
rect 340 -47196 357 -47179
rect 91 -47196 108 -47179
rect 589 -47196 606 -47179
rect 838 -47338 855 -47321
rect 340 -47338 357 -47321
rect 91 -47338 108 -47321
rect 589 -47338 606 -47321
rect 838 -47480 855 -47463
rect 340 -47480 357 -47463
rect 91 -47480 108 -47463
rect 589 -47480 606 -47463
rect 838 -47622 855 -47605
rect 340 -47622 357 -47605
rect 91 -47622 108 -47605
rect 589 -47622 606 -47605
rect 838 -47764 855 -47747
rect 340 -47764 357 -47747
rect 91 -47764 108 -47747
rect 589 -47764 606 -47747
rect 838 -47906 855 -47889
rect 340 -47906 357 -47889
rect 91 -47906 108 -47889
rect 838 -48048 855 -48031
rect 340 -48048 357 -48031
rect 91 -48048 108 -48031
rect 589 -48048 606 -48031
rect 838 -48190 855 -48173
rect 340 -48190 357 -48173
rect 91 -48190 108 -48173
rect 589 -48190 606 -48173
rect 838 -48332 855 -48315
rect 340 -48332 357 -48315
rect 91 -48332 108 -48315
rect 589 -48332 606 -48315
rect 838 -48474 855 -48457
rect 340 -48474 357 -48457
rect 91 -48474 108 -48457
rect 589 -48474 606 -48457
rect 838 -48616 855 -48599
rect 340 -48616 357 -48599
rect 91 -48616 108 -48599
rect 589 -48616 606 -48599
rect 838 -48758 855 -48741
rect 340 -48758 357 -48741
rect 91 -48758 108 -48741
rect 589 -48758 606 -48741
rect 838 -48900 855 -48883
rect 340 -48900 357 -48883
rect 91 -48900 108 -48883
rect 589 -48900 606 -48883
rect 838 -49042 855 -49025
rect 340 -49042 357 -49025
rect 91 -49042 108 -49025
rect 838 -49184 855 -49167
rect 340 -49184 357 -49167
rect 91 -49184 108 -49167
rect 589 -49184 606 -49167
rect 838 -49326 855 -49309
rect 340 -49326 357 -49309
rect 91 -49326 108 -49309
rect 589 -49326 606 -49309
rect 838 -49468 855 -49451
rect 340 -49468 357 -49451
rect 91 -49468 108 -49451
rect 589 -49468 606 -49451
rect 838 -49610 855 -49593
rect 340 -49610 357 -49593
rect 91 -49610 108 -49593
rect 589 -49610 606 -49593
rect 838 -49752 855 -49735
rect 340 -49752 357 -49735
rect 91 -49752 108 -49735
rect 589 -49752 606 -49735
rect 838 -49894 855 -49877
rect 340 -49894 357 -49877
rect 91 -49894 108 -49877
rect 589 -49894 606 -49877
rect 838 -50036 855 -50019
rect 340 -50036 357 -50019
rect 91 -50036 108 -50019
rect 589 -50036 606 -50019
rect 838 -50178 855 -50161
rect 91 -50178 108 -50161
rect 838 -50320 855 -50303
rect 91 -50320 108 -50303
rect 589 -50320 606 -50303
rect 838 -50462 855 -50445
rect 91 -50462 108 -50445
rect 589 -50462 606 -50445
rect 838 -50604 855 -50587
rect 91 -50604 108 -50587
rect 589 -50604 606 -50587
rect 838 -50746 855 -50729
rect 91 -50746 108 -50729
rect 589 -50746 606 -50729
rect 838 -50888 855 -50871
rect 91 -50888 108 -50871
rect 589 -50888 606 -50871
rect 838 -51030 855 -51013
rect 91 -51030 108 -51013
rect 589 -51030 606 -51013
rect 838 -51172 855 -51155
rect 340 -51172 357 -51155
rect 91 -51172 108 -51155
rect 589 -51172 606 -51155
rect 838 -51314 855 -51297
rect 340 -51314 357 -51297
rect 91 -51314 108 -51297
rect 838 -51456 855 -51439
rect 340 -51456 357 -51439
rect 91 -51456 108 -51439
rect 589 -51456 606 -51439
rect 838 -51598 855 -51581
rect 340 -51598 357 -51581
rect 91 -51598 108 -51581
rect 589 -51598 606 -51581
rect 838 -51740 855 -51723
rect 340 -51740 357 -51723
rect 91 -51740 108 -51723
rect 589 -51740 606 -51723
rect 838 -51882 855 -51865
rect 340 -51882 357 -51865
rect 91 -51882 108 -51865
rect 589 -51882 606 -51865
rect 838 -52024 855 -52007
rect 340 -52024 357 -52007
rect 91 -52024 108 -52007
rect 589 -52024 606 -52007
rect 838 -52166 855 -52149
rect 340 -52166 357 -52149
rect 91 -52166 108 -52149
rect 589 -52166 606 -52149
rect 838 -52308 855 -52291
rect 340 -52308 357 -52291
rect 91 -52308 108 -52291
rect 589 -52308 606 -52291
rect 838 -52450 855 -52433
rect 340 -52450 357 -52433
rect 91 -52450 108 -52433
rect 838 -52592 855 -52575
rect 340 -52592 357 -52575
rect 91 -52592 108 -52575
rect 589 -52592 606 -52575
rect 838 -52734 855 -52717
rect 340 -52734 357 -52717
rect 91 -52734 108 -52717
rect 589 -52734 606 -52717
rect 838 -52876 855 -52859
rect 340 -52876 357 -52859
rect 91 -52876 108 -52859
rect 589 -52876 606 -52859
rect 838 -53018 855 -53001
rect 340 -53018 357 -53001
rect 91 -53018 108 -53001
rect 589 -53018 606 -53001
rect 838 -53160 855 -53143
rect 340 -53160 357 -53143
rect 91 -53160 108 -53143
rect 589 -53160 606 -53143
rect 838 -53302 855 -53285
rect 340 -53302 357 -53285
rect 91 -53302 108 -53285
rect 589 -53302 606 -53285
rect 838 -53444 855 -53427
rect 340 -53444 357 -53427
rect 91 -53444 108 -53427
rect 589 -53444 606 -53427
rect 838 -53586 855 -53569
rect 340 -53586 357 -53569
rect 91 -53586 108 -53569
rect 838 -53728 855 -53711
rect 340 -53728 357 -53711
rect 91 -53728 108 -53711
rect 589 -53728 606 -53711
rect 838 -53870 855 -53853
rect 340 -53870 357 -53853
rect 91 -53870 108 -53853
rect 589 -53870 606 -53853
rect 838 -54012 855 -53995
rect 340 -54012 357 -53995
rect 91 -54012 108 -53995
rect 589 -54012 606 -53995
rect 838 -54154 855 -54137
rect 340 -54154 357 -54137
rect 91 -54154 108 -54137
rect 589 -54154 606 -54137
rect 838 -54296 855 -54279
rect 340 -54296 357 -54279
rect 91 -54296 108 -54279
rect 589 -54296 606 -54279
rect 838 -54438 855 -54421
rect 340 -54438 357 -54421
rect 91 -54438 108 -54421
rect 589 -54438 606 -54421
rect 838 -54864 855 -54847
rect 838 -55006 855 -54989
rect 838 -55148 855 -55131
rect 589 -55290 606 -55273
rect 838 -55290 855 -55273
rect 838 -55432 855 -55415
rect 589 -55432 606 -55415
rect 838 -55574 855 -55557
rect 589 -55574 606 -55557
rect 838 -55716 855 -55699
rect 589 -55716 606 -55699
rect 838 -55858 855 -55841
rect 589 -55858 606 -55841
rect 838 -56000 855 -55983
rect 340 -56000 357 -55983
rect 589 -56000 606 -55983
rect 838 -56142 855 -56125
rect 340 -56142 357 -56125
rect 589 -56142 606 -56125
rect 838 -56284 855 -56267
rect 340 -56284 357 -56267
rect 589 -56284 606 -56267
rect 838 -56426 855 -56409
rect 340 -56426 357 -56409
rect 589 -56426 606 -56409
rect 838 -56568 855 -56551
rect 340 -56568 357 -56551
rect 589 -56568 606 -56551
rect 838 -56710 855 -56693
rect 340 -56710 357 -56693
rect 838 -56852 855 -56835
rect 340 -56852 357 -56835
rect 589 -56852 606 -56835
rect 838 -56994 855 -56977
rect 340 -56994 357 -56977
rect 589 -56994 606 -56977
rect 838 -57136 855 -57119
rect 340 -57136 357 -57119
rect 589 -57136 606 -57119
rect 838 -57278 855 -57261
rect 340 -57278 357 -57261
rect 589 -57278 606 -57261
rect 838 -57420 855 -57403
rect 340 -57420 357 -57403
rect 589 -57420 606 -57403
rect 838 -57562 855 -57545
rect 340 -57562 357 -57545
rect 91 -57562 108 -57545
rect 589 -57562 606 -57545
rect 838 -57704 855 -57687
rect 91 -57704 108 -57687
rect 589 -57704 606 -57687
rect 838 -57846 855 -57829
rect 91 -57846 108 -57829
rect 589 -57846 606 -57829
rect 838 -57988 855 -57971
rect 340 -57988 357 -57971
rect 91 -57988 108 -57971
rect 589 -57988 606 -57971
rect 838 -58130 855 -58113
rect 340 -58130 357 -58113
rect 91 -58130 108 -58113
rect 589 -58130 606 -58113
rect 838 -58272 855 -58255
rect 340 -58272 357 -58255
rect 91 -58272 108 -58255
rect 589 -58272 606 -58255
rect 838 -58414 855 -58397
rect 340 -58414 357 -58397
rect 91 -58414 108 -58397
rect 589 -58414 606 -58397
rect 838 -58556 855 -58539
rect 340 -58556 357 -58539
rect 91 -58556 108 -58539
rect 589 -58556 606 -58539
rect 838 -58698 855 -58681
rect 340 -58698 357 -58681
rect 91 -58698 108 -58681
rect 589 -58698 606 -58681
rect 838 -58840 855 -58823
rect 340 -58840 357 -58823
rect 91 -58840 108 -58823
rect 589 -58840 606 -58823
rect 838 -58982 855 -58965
rect 340 -58982 357 -58965
rect 91 -58982 108 -58965
rect 589 -58982 606 -58965
rect 838 -59124 855 -59107
rect 91 -59124 108 -59107
rect 838 -59266 855 -59249
rect 91 -59266 108 -59249
rect 589 -59266 606 -59249
rect 838 -59408 855 -59391
rect 91 -59408 108 -59391
rect 589 -59408 606 -59391
rect 838 -59550 855 -59533
rect 340 -59550 357 -59533
rect 91 -59550 108 -59533
rect 589 -59550 606 -59533
rect 838 -59692 855 -59675
rect 340 -59692 357 -59675
rect 91 -59692 108 -59675
rect 589 -59692 606 -59675
rect 838 -59834 855 -59817
rect 340 -59834 357 -59817
rect 91 -59834 108 -59817
rect 589 -59834 606 -59817
rect 838 -59976 855 -59959
rect 340 -59976 357 -59959
rect 91 -59976 108 -59959
rect 589 -59976 606 -59959
rect 838 -60118 855 -60101
rect 340 -60118 357 -60101
rect 91 -60118 108 -60101
rect 589 -60118 606 -60101
rect 838 -60260 855 -60243
rect 340 -60260 357 -60243
rect 91 -60260 108 -60243
rect 838 -60402 855 -60385
rect 340 -60402 357 -60385
rect 91 -60402 108 -60385
rect 589 -60402 606 -60385
rect 838 -60544 855 -60527
rect 340 -60544 357 -60527
rect 91 -60544 108 -60527
rect 589 -60544 606 -60527
rect 838 -60686 855 -60669
rect 91 -60686 108 -60669
rect 589 -60686 606 -60669
rect 838 -60828 855 -60811
rect 91 -60828 108 -60811
rect 589 -60828 606 -60811
rect 838 -60970 855 -60953
rect 91 -60970 108 -60953
rect 589 -60970 606 -60953
rect 838 -61112 855 -61095
rect 340 -61112 357 -61095
rect 91 -61112 108 -61095
rect 838 -61254 855 -61237
rect 340 -61254 357 -61237
rect 91 -61254 108 -61237
rect 589 -61254 606 -61237
rect 838 -61396 855 -61379
rect 340 -61396 357 -61379
rect 91 -61396 108 -61379
rect 589 -61396 606 -61379
rect 838 -61538 855 -61521
rect 340 -61538 357 -61521
rect 91 -61538 108 -61521
rect 589 -61538 606 -61521
rect 838 -61680 855 -61663
rect 340 -61680 357 -61663
rect 91 -61680 108 -61663
rect 589 -61680 606 -61663
rect 838 -61822 855 -61805
rect 340 -61822 357 -61805
rect 91 -61822 108 -61805
rect 589 -61822 606 -61805
rect 838 -61964 855 -61947
rect 340 -61964 357 -61947
rect 91 -61964 108 -61947
rect 589 -61964 606 -61947
rect 838 -62106 855 -62089
rect 340 -62106 357 -62089
rect 91 -62106 108 -62089
rect 589 -62106 606 -62089
rect 838 -62248 855 -62231
rect 340 -62248 357 -62231
rect 91 -62248 108 -62231
rect 838 -62390 855 -62373
rect 340 -62390 357 -62373
rect 91 -62390 108 -62373
rect 589 -62390 606 -62373
rect 838 -62532 855 -62515
rect 340 -62532 357 -62515
rect 91 -62532 108 -62515
rect 589 -62532 606 -62515
rect 838 -62674 855 -62657
rect 340 -62674 357 -62657
rect 91 -62674 108 -62657
rect 589 -62674 606 -62657
rect 838 -62816 855 -62799
rect 340 -62816 357 -62799
rect 91 -62816 108 -62799
rect 589 -62816 606 -62799
rect 838 -62958 855 -62941
rect 340 -62958 357 -62941
rect 91 -62958 108 -62941
rect 589 -62958 606 -62941
rect 838 -63100 855 -63083
rect 340 -63100 357 -63083
rect 91 -63100 108 -63083
rect 589 -63100 606 -63083
rect 838 -63242 855 -63225
rect 340 -63242 357 -63225
rect 91 -63242 108 -63225
rect 589 -63242 606 -63225
rect 838 -63384 855 -63367
rect 340 -63384 357 -63367
rect 91 -63384 108 -63367
rect 589 -63384 606 -63367
rect 838 -63526 855 -63509
rect 340 -63526 357 -63509
rect 91 -63526 108 -63509
rect 589 -63526 606 -63509
rect 838 -63668 855 -63651
rect 340 -63668 357 -63651
rect 91 -63668 108 -63651
rect 589 -63668 606 -63651
rect 838 -63810 855 -63793
rect 340 -63810 357 -63793
rect 91 -63810 108 -63793
rect 589 -63810 606 -63793
rect 838 -63952 855 -63935
rect 340 -63952 357 -63935
rect 91 -63952 108 -63935
rect 589 -63952 606 -63935
rect 838 -64094 855 -64077
rect 340 -64094 357 -64077
rect 91 -64094 108 -64077
rect 589 -64094 606 -64077
rect 838 -64236 855 -64219
rect 340 -64236 357 -64219
rect 91 -64236 108 -64219
rect 589 -64236 606 -64219
rect 838 -64378 855 -64361
rect 340 -64378 357 -64361
rect 91 -64378 108 -64361
rect 589 -64378 606 -64361
rect 838 -64520 855 -64503
rect 340 -64520 357 -64503
rect 91 -64520 108 -64503
rect 589 -64520 606 -64503
rect 838 -64662 855 -64645
rect 340 -64662 357 -64645
rect 91 -64662 108 -64645
rect 589 -64662 606 -64645
rect 838 -64804 855 -64787
rect 340 -64804 357 -64787
rect 91 -64804 108 -64787
rect 589 -64804 606 -64787
rect 838 -64946 855 -64929
rect 340 -64946 357 -64929
rect 91 -64946 108 -64929
rect 838 -65088 855 -65071
rect 340 -65088 357 -65071
rect 91 -65088 108 -65071
rect 589 -65088 606 -65071
rect 838 -65230 855 -65213
rect 340 -65230 357 -65213
rect 91 -65230 108 -65213
rect 589 -65230 606 -65213
rect 838 -65372 855 -65355
rect 340 -65372 357 -65355
rect 91 -65372 108 -65355
rect 589 -65372 606 -65355
rect 838 -65514 855 -65497
rect 340 -65514 357 -65497
rect 91 -65514 108 -65497
rect 589 -65514 606 -65497
rect 838 -65656 855 -65639
rect 340 -65656 357 -65639
rect 91 -65656 108 -65639
rect 838 -65798 855 -65781
rect 340 -65798 357 -65781
rect 91 -65798 108 -65781
rect 589 -65798 606 -65781
rect 838 -65940 855 -65923
rect 340 -65940 357 -65923
rect 91 -65940 108 -65923
rect 589 -65940 606 -65923
rect 838 -66082 855 -66065
rect 340 -66082 357 -66065
rect 91 -66082 108 -66065
rect 589 -66082 606 -66065
rect 838 -66224 855 -66207
rect 340 -66224 357 -66207
rect 91 -66224 108 -66207
rect 589 -66224 606 -66207
rect 838 -66366 855 -66349
rect 91 -66366 108 -66349
rect 589 -66366 606 -66349
rect 838 -66508 855 -66491
rect 91 -66508 108 -66491
rect 589 -66508 606 -66491
rect 838 -66650 855 -66633
rect 340 -66650 357 -66633
rect 91 -66650 108 -66633
rect 589 -66650 606 -66633
rect 838 -66792 855 -66775
rect 340 -66792 357 -66775
rect 91 -66792 108 -66775
rect 589 -66792 606 -66775
rect 838 -66934 855 -66917
rect 340 -66934 357 -66917
rect 91 -66934 108 -66917
rect 589 -66934 606 -66917
rect 838 -67076 855 -67059
rect 340 -67076 357 -67059
rect 91 -67076 108 -67059
rect 589 -67076 606 -67059
rect 838 -67218 855 -67201
rect 340 -67218 357 -67201
rect 91 -67218 108 -67201
rect 589 -67218 606 -67201
rect 838 -67360 855 -67343
rect 340 -67360 357 -67343
rect 91 -67360 108 -67343
rect 589 -67360 606 -67343
rect 838 -67502 855 -67485
rect 340 -67502 357 -67485
rect 91 -67502 108 -67485
rect 589 -67502 606 -67485
rect 838 -67644 855 -67627
rect 340 -67644 357 -67627
rect 91 -67644 108 -67627
rect 589 -67644 606 -67627
rect 838 -67786 855 -67769
rect 340 -67786 357 -67769
rect 91 -67786 108 -67769
rect 589 -67786 606 -67769
rect 838 -67928 855 -67911
rect 91 -67928 108 -67911
rect 589 -67928 606 -67911
rect 838 -68070 855 -68053
rect 91 -68070 108 -68053
rect 589 -68070 606 -68053
rect 340 -68212 357 -68195
rect 91 -68212 108 -68195
rect 589 -68212 606 -68195
rect 838 -68354 855 -68337
rect 340 -68354 357 -68337
rect 91 -68354 108 -68337
rect 589 -68354 606 -68337
rect 838 -68496 855 -68479
rect 340 -68496 357 -68479
rect 91 -68496 108 -68479
rect 838 -68638 855 -68621
rect 340 -68638 357 -68621
rect 91 -68638 108 -68621
rect 589 -68638 606 -68621
rect 838 -68780 855 -68763
rect 340 -68780 357 -68763
rect 91 -68780 108 -68763
rect 589 -68780 606 -68763
rect 838 -68922 855 -68905
rect 340 -68922 357 -68905
rect 91 -68922 108 -68905
rect 589 -68922 606 -68905
rect 838 -69064 855 -69047
rect 340 -69064 357 -69047
rect 91 -69064 108 -69047
rect 589 -69064 606 -69047
rect 838 -69206 855 -69189
rect 340 -69206 357 -69189
rect 91 -69206 108 -69189
rect 589 -69206 606 -69189
rect 838 -69348 855 -69331
rect 91 -69348 108 -69331
rect 589 -69348 606 -69331
rect 838 -69490 855 -69473
rect 91 -69490 108 -69473
rect 589 -69490 606 -69473
rect 838 -69632 855 -69615
rect 91 -69632 108 -69615
rect 838 -69774 855 -69757
rect 340 -69774 357 -69757
rect 589 -69774 606 -69757
rect 838 -69916 855 -69899
rect 340 -69916 357 -69899
rect 589 -69916 606 -69899
rect 838 -70058 855 -70041
rect 340 -70058 357 -70041
rect 589 -70058 606 -70041
rect 838 -70200 855 -70183
rect 340 -70200 357 -70183
rect 589 -70200 606 -70183
rect 838 -70342 855 -70325
rect 340 -70342 357 -70325
rect 589 -70342 606 -70325
rect 838 -70484 855 -70467
rect 340 -70484 357 -70467
rect 589 -70484 606 -70467
rect 838 -70626 855 -70609
rect 340 -70626 357 -70609
rect 589 -70626 606 -70609
rect 838 -70768 855 -70751
rect 340 -70768 357 -70751
rect 589 -70768 606 -70751
rect 838 -70910 855 -70893
rect 340 -70910 357 -70893
rect 589 -70910 606 -70893
rect 838 -71052 855 -71035
rect 340 -71052 357 -71035
rect 589 -71052 606 -71035
rect 838 -71194 855 -71177
rect 340 -71194 357 -71177
rect 838 -71336 855 -71319
rect 589 -71336 606 -71319
rect 838 -71478 855 -71461
rect 589 -71478 606 -71461
rect 838 -71620 855 -71603
rect 589 -71620 606 -71603
rect 838 -71762 855 -71745
rect 589 -71762 606 -71745
rect 589 -71904 606 -71887
rect 838 -71904 855 -71887
rect 838 -72046 855 -72029
rect 589 -72046 606 -72029
rect 838 -72188 855 -72171
rect 838 -72330 855 -72313
rect 838 -72472 855 -72455
rect 921 -9069 938 -9052
rect 8 -9069 25 -9052
rect 672 -9069 689 -9052
rect 506 -9069 523 -9052
rect 423 -9069 440 -9052
rect 257 -9069 274 -9052
rect 174 -9069 191 -9052
rect 755 -9069 772 -9052
rect 921 -9211 938 -9194
rect 8 -9211 25 -9194
rect 672 -9211 689 -9194
rect 506 -9211 523 -9194
rect 423 -9211 440 -9194
rect 257 -9211 274 -9194
rect 174 -9211 191 -9194
rect 755 -9211 772 -9194
rect 921 -9353 938 -9336
rect 8 -9353 25 -9336
rect 672 -9353 689 -9336
rect 506 -9353 523 -9336
rect 423 -9353 440 -9336
rect 257 -9353 274 -9336
rect 174 -9353 191 -9336
rect 755 -9353 772 -9336
rect 921 -9495 938 -9478
rect 8 -9495 25 -9478
rect 672 -9495 689 -9478
rect 506 -9495 523 -9478
rect 423 -9495 440 -9478
rect 257 -9495 274 -9478
rect 174 -9495 191 -9478
rect 755 -9495 772 -9478
rect 921 -9637 938 -9620
rect 8 -9637 25 -9620
rect 672 -9637 689 -9620
rect 506 -9637 523 -9620
rect 423 -9637 440 -9620
rect 257 -9637 274 -9620
rect 174 -9637 191 -9620
rect 755 -9637 772 -9620
rect 921 -9779 938 -9762
rect 8 -9779 25 -9762
rect 672 -9779 689 -9762
rect 506 -9779 523 -9762
rect 423 -9779 440 -9762
rect 257 -9779 274 -9762
rect 174 -9779 191 -9762
rect 755 -9779 772 -9762
rect 921 -9921 938 -9904
rect 8 -9921 25 -9904
rect 672 -9921 689 -9904
rect 506 -9921 523 -9904
rect 423 -9921 440 -9904
rect 257 -9921 274 -9904
rect 174 -9921 191 -9904
rect 755 -9921 772 -9904
rect 921 -10063 938 -10046
rect 8 -10063 25 -10046
rect 672 -10063 689 -10046
rect 506 -10063 523 -10046
rect 423 -10063 440 -10046
rect 257 -10063 274 -10046
rect 174 -10063 191 -10046
rect 755 -10063 772 -10046
rect 921 -10205 938 -10188
rect 8 -10205 25 -10188
rect 672 -10205 689 -10188
rect 506 -10205 523 -10188
rect 423 -10205 440 -10188
rect 257 -10205 274 -10188
rect 174 -10205 191 -10188
rect 755 -10205 772 -10188
rect 921 -10347 938 -10330
rect 8 -10347 25 -10330
rect 672 -10347 689 -10330
rect 506 -10347 523 -10330
rect 423 -10347 440 -10330
rect 257 -10347 274 -10330
rect 174 -10347 191 -10330
rect 755 -10347 772 -10330
rect 921 -10489 938 -10472
rect 8 -10489 25 -10472
rect 672 -10489 689 -10472
rect 506 -10489 523 -10472
rect 423 -10489 440 -10472
rect 257 -10489 274 -10472
rect 174 -10489 191 -10472
rect 755 -10489 772 -10472
rect 921 -10631 938 -10614
rect 8 -10631 25 -10614
rect 672 -10631 689 -10614
rect 506 -10631 523 -10614
rect 423 -10631 440 -10614
rect 257 -10631 274 -10614
rect 174 -10631 191 -10614
rect 755 -10631 772 -10614
rect 921 -10773 938 -10756
rect 8 -10773 25 -10756
rect 672 -10773 689 -10756
rect 506 -10773 523 -10756
rect 423 -10773 440 -10756
rect 257 -10773 274 -10756
rect 174 -10773 191 -10756
rect 755 -10773 772 -10756
rect 921 -10915 938 -10898
rect 8 -10915 25 -10898
rect 672 -10915 689 -10898
rect 506 -10915 523 -10898
rect 423 -10915 440 -10898
rect 257 -10915 274 -10898
rect 174 -10915 191 -10898
rect 755 -10915 772 -10898
rect 921 -11057 938 -11040
rect 8 -11057 25 -11040
rect 672 -11057 689 -11040
rect 506 -11057 523 -11040
rect 423 -11057 440 -11040
rect 257 -11057 274 -11040
rect 174 -11057 191 -11040
rect 755 -11057 772 -11040
rect 921 -11199 938 -11182
rect 8 -11199 25 -11182
rect 672 -11199 689 -11182
rect 506 -11199 523 -11182
rect 423 -11199 440 -11182
rect 257 -11199 274 -11182
rect 174 -11199 191 -11182
rect 755 -11199 772 -11182
rect 921 -11341 938 -11324
rect 8 -11341 25 -11324
rect 672 -11341 689 -11324
rect 506 -11341 523 -11324
rect 423 -11341 440 -11324
rect 257 -11341 274 -11324
rect 174 -11341 191 -11324
rect 755 -11341 772 -11324
rect 921 -11483 938 -11466
rect 8 -11483 25 -11466
rect 672 -11483 689 -11466
rect 506 -11483 523 -11466
rect 423 -11483 440 -11466
rect 257 -11483 274 -11466
rect 174 -11483 191 -11466
rect 755 -11483 772 -11466
rect 921 -11625 938 -11608
rect 8 -11625 25 -11608
rect 672 -11625 689 -11608
rect 506 -11625 523 -11608
rect 423 -11625 440 -11608
rect 257 -11625 274 -11608
rect 174 -11625 191 -11608
rect 755 -11625 772 -11608
rect 921 -11767 938 -11750
rect 8 -11767 25 -11750
rect 672 -11767 689 -11750
rect 506 -11767 523 -11750
rect 423 -11767 440 -11750
rect 257 -11767 274 -11750
rect 174 -11767 191 -11750
rect 755 -11767 772 -11750
rect 921 -11909 938 -11892
rect 8 -11909 25 -11892
rect 672 -11909 689 -11892
rect 506 -11909 523 -11892
rect 423 -11909 440 -11892
rect 257 -11909 274 -11892
rect 174 -11909 191 -11892
rect 755 -11909 772 -11892
rect 921 -12051 938 -12034
rect 8 -12051 25 -12034
rect 672 -12051 689 -12034
rect 506 -12051 523 -12034
rect 423 -12051 440 -12034
rect 257 -12051 274 -12034
rect 174 -12051 191 -12034
rect 755 -12051 772 -12034
rect 921 -12193 938 -12176
rect 8 -12193 25 -12176
rect 672 -12193 689 -12176
rect 506 -12193 523 -12176
rect 423 -12193 440 -12176
rect 257 -12193 274 -12176
rect 174 -12193 191 -12176
rect 755 -12193 772 -12176
rect 921 -12335 938 -12318
rect 8 -12335 25 -12318
rect 672 -12335 689 -12318
rect 506 -12335 523 -12318
rect 423 -12335 440 -12318
rect 257 -12335 274 -12318
rect 174 -12335 191 -12318
rect 755 -12335 772 -12318
rect 921 -12477 938 -12460
rect 8 -12477 25 -12460
rect 672 -12477 689 -12460
rect 506 -12477 523 -12460
rect 423 -12477 440 -12460
rect 257 -12477 274 -12460
rect 174 -12477 191 -12460
rect 755 -12477 772 -12460
rect 921 -12619 938 -12602
rect 8 -12619 25 -12602
rect 672 -12619 689 -12602
rect 506 -12619 523 -12602
rect 423 -12619 440 -12602
rect 257 -12619 274 -12602
rect 174 -12619 191 -12602
rect 755 -12619 772 -12602
rect 921 -12761 938 -12744
rect 8 -12761 25 -12744
rect 672 -12761 689 -12744
rect 506 -12761 523 -12744
rect 423 -12761 440 -12744
rect 257 -12761 274 -12744
rect 174 -12761 191 -12744
rect 755 -12761 772 -12744
rect 921 -12903 938 -12886
rect 8 -12903 25 -12886
rect 672 -12903 689 -12886
rect 506 -12903 523 -12886
rect 423 -12903 440 -12886
rect 257 -12903 274 -12886
rect 174 -12903 191 -12886
rect 755 -12903 772 -12886
rect 921 -13045 938 -13028
rect 8 -13045 25 -13028
rect 672 -13045 689 -13028
rect 506 -13045 523 -13028
rect 423 -13045 440 -13028
rect 257 -13045 274 -13028
rect 174 -13045 191 -13028
rect 755 -13045 772 -13028
rect 921 -13187 938 -13170
rect 8 -13187 25 -13170
rect 672 -13187 689 -13170
rect 506 -13187 523 -13170
rect 423 -13187 440 -13170
rect 257 -13187 274 -13170
rect 174 -13187 191 -13170
rect 755 -13187 772 -13170
rect 921 -13329 938 -13312
rect 8 -13329 25 -13312
rect 672 -13329 689 -13312
rect 506 -13329 523 -13312
rect 423 -13329 440 -13312
rect 257 -13329 274 -13312
rect 174 -13329 191 -13312
rect 755 -13329 772 -13312
rect 921 -13471 938 -13454
rect 8 -13471 25 -13454
rect 672 -13471 689 -13454
rect 506 -13471 523 -13454
rect 423 -13471 440 -13454
rect 257 -13471 274 -13454
rect 174 -13471 191 -13454
rect 755 -13471 772 -13454
rect 921 -13613 938 -13596
rect 8 -13613 25 -13596
rect 672 -13613 689 -13596
rect 506 -13613 523 -13596
rect 423 -13613 440 -13596
rect 257 -13613 274 -13596
rect 174 -13613 191 -13596
rect 755 -13613 772 -13596
rect 921 -13755 938 -13738
rect 8 -13755 25 -13738
rect 672 -13755 689 -13738
rect 506 -13755 523 -13738
rect 423 -13755 440 -13738
rect 257 -13755 274 -13738
rect 174 -13755 191 -13738
rect 755 -13755 772 -13738
rect 921 -13897 938 -13880
rect 8 -13897 25 -13880
rect 672 -13897 689 -13880
rect 506 -13897 523 -13880
rect 423 -13897 440 -13880
rect 257 -13897 274 -13880
rect 174 -13897 191 -13880
rect 755 -13897 772 -13880
rect 921 -14039 938 -14022
rect 8 -14039 25 -14022
rect 672 -14039 689 -14022
rect 506 -14039 523 -14022
rect 423 -14039 440 -14022
rect 257 -14039 274 -14022
rect 174 -14039 191 -14022
rect 755 -14039 772 -14022
rect 921 -14181 938 -14164
rect 8 -14181 25 -14164
rect 672 -14181 689 -14164
rect 506 -14181 523 -14164
rect 423 -14181 440 -14164
rect 257 -14181 274 -14164
rect 174 -14181 191 -14164
rect 755 -14181 772 -14164
rect 921 -14323 938 -14306
rect 8 -14323 25 -14306
rect 672 -14323 689 -14306
rect 506 -14323 523 -14306
rect 423 -14323 440 -14306
rect 257 -14323 274 -14306
rect 174 -14323 191 -14306
rect 755 -14323 772 -14306
rect 921 -14465 938 -14448
rect 8 -14465 25 -14448
rect 672 -14465 689 -14448
rect 506 -14465 523 -14448
rect 423 -14465 440 -14448
rect 257 -14465 274 -14448
rect 174 -14465 191 -14448
rect 755 -14465 772 -14448
rect 921 -14607 938 -14590
rect 8 -14607 25 -14590
rect 672 -14607 689 -14590
rect 506 -14607 523 -14590
rect 423 -14607 440 -14590
rect 257 -14607 274 -14590
rect 174 -14607 191 -14590
rect 755 -14607 772 -14590
rect 921 -14749 938 -14732
rect 8 -14749 25 -14732
rect 672 -14749 689 -14732
rect 506 -14749 523 -14732
rect 423 -14749 440 -14732
rect 257 -14749 274 -14732
rect 174 -14749 191 -14732
rect 755 -14749 772 -14732
rect 921 -14891 938 -14874
rect 8 -14891 25 -14874
rect 672 -14891 689 -14874
rect 506 -14891 523 -14874
rect 423 -14891 440 -14874
rect 257 -14891 274 -14874
rect 174 -14891 191 -14874
rect 755 -14891 772 -14874
rect 921 -15033 938 -15016
rect 8 -15033 25 -15016
rect 672 -15033 689 -15016
rect 506 -15033 523 -15016
rect 423 -15033 440 -15016
rect 257 -15033 274 -15016
rect 174 -15033 191 -15016
rect 755 -15033 772 -15016
rect 921 -15175 938 -15158
rect 8 -15175 25 -15158
rect 672 -15175 689 -15158
rect 506 -15175 523 -15158
rect 423 -15175 440 -15158
rect 257 -15175 274 -15158
rect 174 -15175 191 -15158
rect 755 -15175 772 -15158
rect 921 -15317 938 -15300
rect 8 -15317 25 -15300
rect 672 -15317 689 -15300
rect 506 -15317 523 -15300
rect 423 -15317 440 -15300
rect 257 -15317 274 -15300
rect 174 -15317 191 -15300
rect 755 -15317 772 -15300
rect 921 -15459 938 -15442
rect 8 -15459 25 -15442
rect 672 -15459 689 -15442
rect 506 -15459 523 -15442
rect 423 -15459 440 -15442
rect 257 -15459 274 -15442
rect 174 -15459 191 -15442
rect 755 -15459 772 -15442
rect 921 -15601 938 -15584
rect 8 -15601 25 -15584
rect 672 -15601 689 -15584
rect 506 -15601 523 -15584
rect 423 -15601 440 -15584
rect 257 -15601 274 -15584
rect 174 -15601 191 -15584
rect 755 -15601 772 -15584
rect 921 -15743 938 -15726
rect 8 -15743 25 -15726
rect 672 -15743 689 -15726
rect 506 -15743 523 -15726
rect 423 -15743 440 -15726
rect 257 -15743 274 -15726
rect 174 -15743 191 -15726
rect 755 -15743 772 -15726
rect 921 -15885 938 -15868
rect 8 -15885 25 -15868
rect 672 -15885 689 -15868
rect 506 -15885 523 -15868
rect 423 -15885 440 -15868
rect 257 -15885 274 -15868
rect 174 -15885 191 -15868
rect 755 -15885 772 -15868
rect 921 -16027 938 -16010
rect 8 -16027 25 -16010
rect 672 -16027 689 -16010
rect 506 -16027 523 -16010
rect 423 -16027 440 -16010
rect 257 -16027 274 -16010
rect 174 -16027 191 -16010
rect 755 -16027 772 -16010
rect 921 -16169 938 -16152
rect 8 -16169 25 -16152
rect 672 -16169 689 -16152
rect 506 -16169 523 -16152
rect 423 -16169 440 -16152
rect 257 -16169 274 -16152
rect 174 -16169 191 -16152
rect 755 -16169 772 -16152
rect 921 -16311 938 -16294
rect 8 -16311 25 -16294
rect 672 -16311 689 -16294
rect 506 -16311 523 -16294
rect 423 -16311 440 -16294
rect 257 -16311 274 -16294
rect 174 -16311 191 -16294
rect 755 -16311 772 -16294
rect 921 -16453 938 -16436
rect 8 -16453 25 -16436
rect 672 -16453 689 -16436
rect 506 -16453 523 -16436
rect 423 -16453 440 -16436
rect 257 -16453 274 -16436
rect 174 -16453 191 -16436
rect 755 -16453 772 -16436
rect 921 -16595 938 -16578
rect 8 -16595 25 -16578
rect 672 -16595 689 -16578
rect 506 -16595 523 -16578
rect 423 -16595 440 -16578
rect 257 -16595 274 -16578
rect 174 -16595 191 -16578
rect 755 -16595 772 -16578
rect 921 -16737 938 -16720
rect 8 -16737 25 -16720
rect 672 -16737 689 -16720
rect 506 -16737 523 -16720
rect 423 -16737 440 -16720
rect 257 -16737 274 -16720
rect 174 -16737 191 -16720
rect 755 -16737 772 -16720
rect 921 -16879 938 -16862
rect 8 -16879 25 -16862
rect 672 -16879 689 -16862
rect 506 -16879 523 -16862
rect 423 -16879 440 -16862
rect 257 -16879 274 -16862
rect 174 -16879 191 -16862
rect 755 -16879 772 -16862
rect 921 -17021 938 -17004
rect 8 -17021 25 -17004
rect 672 -17021 689 -17004
rect 506 -17021 523 -17004
rect 423 -17021 440 -17004
rect 257 -17021 274 -17004
rect 174 -17021 191 -17004
rect 755 -17021 772 -17004
rect 921 -17163 938 -17146
rect 8 -17163 25 -17146
rect 672 -17163 689 -17146
rect 506 -17163 523 -17146
rect 423 -17163 440 -17146
rect 257 -17163 274 -17146
rect 174 -17163 191 -17146
rect 755 -17163 772 -17146
rect 921 -17305 938 -17288
rect 8 -17305 25 -17288
rect 672 -17305 689 -17288
rect 506 -17305 523 -17288
rect 423 -17305 440 -17288
rect 257 -17305 274 -17288
rect 174 -17305 191 -17288
rect 755 -17305 772 -17288
rect 921 -17447 938 -17430
rect 8 -17447 25 -17430
rect 672 -17447 689 -17430
rect 506 -17447 523 -17430
rect 423 -17447 440 -17430
rect 257 -17447 274 -17430
rect 174 -17447 191 -17430
rect 755 -17447 772 -17430
rect 921 -17589 938 -17572
rect 8 -17589 25 -17572
rect 672 -17589 689 -17572
rect 506 -17589 523 -17572
rect 423 -17589 440 -17572
rect 257 -17589 274 -17572
rect 174 -17589 191 -17572
rect 755 -17589 772 -17572
rect 921 -17731 938 -17714
rect 8 -17731 25 -17714
rect 672 -17731 689 -17714
rect 506 -17731 523 -17714
rect 423 -17731 440 -17714
rect 257 -17731 274 -17714
rect 174 -17731 191 -17714
rect 755 -17731 772 -17714
rect 921 -17873 938 -17856
rect 8 -17873 25 -17856
rect 672 -17873 689 -17856
rect 506 -17873 523 -17856
rect 423 -17873 440 -17856
rect 257 -17873 274 -17856
rect 174 -17873 191 -17856
rect 755 -17873 772 -17856
rect 921 -18015 938 -17998
rect 8 -18015 25 -17998
rect 672 -18015 689 -17998
rect 506 -18015 523 -17998
rect 423 -18015 440 -17998
rect 257 -18015 274 -17998
rect 174 -18015 191 -17998
rect 755 -18015 772 -17998
rect 921 -18157 938 -18140
rect 8 -18157 25 -18140
rect 672 -18157 689 -18140
rect 506 -18157 523 -18140
rect 423 -18157 440 -18140
rect 257 -18157 274 -18140
rect 174 -18157 191 -18140
rect 755 -18157 772 -18140
rect 755 -18299 772 -18282
rect 921 -18299 938 -18282
rect 921 -18441 938 -18424
rect 672 -18441 689 -18424
rect 755 -18441 772 -18424
rect 921 -18583 938 -18566
rect 506 -18583 523 -18566
rect 755 -18583 772 -18566
rect 921 -18725 938 -18708
rect 672 -18725 689 -18708
rect 506 -18725 523 -18708
rect 755 -18725 772 -18708
rect 921 -18867 938 -18850
rect 423 -18867 440 -18850
rect 755 -18867 772 -18850
rect 921 -19009 938 -18992
rect 423 -19009 440 -18992
rect 672 -19009 689 -18992
rect 755 -19009 772 -18992
rect 921 -19151 938 -19134
rect 423 -19151 440 -19134
rect 506 -19151 523 -19134
rect 755 -19151 772 -19134
rect 921 -19293 938 -19276
rect 672 -19293 689 -19276
rect 506 -19293 523 -19276
rect 423 -19293 440 -19276
rect 755 -19293 772 -19276
rect 921 -19435 938 -19418
rect 257 -19435 274 -19418
rect 755 -19435 772 -19418
rect 921 -19577 938 -19560
rect 672 -19577 689 -19560
rect 257 -19577 274 -19560
rect 755 -19577 772 -19560
rect 921 -19719 938 -19702
rect 506 -19719 523 -19702
rect 257 -19719 274 -19702
rect 755 -19719 772 -19702
rect 921 -19861 938 -19844
rect 672 -19861 689 -19844
rect 506 -19861 523 -19844
rect 257 -19861 274 -19844
rect 755 -19861 772 -19844
rect 921 -20003 938 -19986
rect 423 -20003 440 -19986
rect 257 -20003 274 -19986
rect 755 -20003 772 -19986
rect 921 -20145 938 -20128
rect 423 -20145 440 -20128
rect 672 -20145 689 -20128
rect 257 -20145 274 -20128
rect 755 -20145 772 -20128
rect 921 -20287 938 -20270
rect 423 -20287 440 -20270
rect 506 -20287 523 -20270
rect 257 -20287 274 -20270
rect 755 -20287 772 -20270
rect 921 -20429 938 -20412
rect 672 -20429 689 -20412
rect 506 -20429 523 -20412
rect 423 -20429 440 -20412
rect 257 -20429 274 -20412
rect 755 -20429 772 -20412
rect 921 -20571 938 -20554
rect 174 -20571 191 -20554
rect 755 -20571 772 -20554
rect 921 -20713 938 -20696
rect 672 -20713 689 -20696
rect 174 -20713 191 -20696
rect 755 -20713 772 -20696
rect 921 -20855 938 -20838
rect 506 -20855 523 -20838
rect 174 -20855 191 -20838
rect 755 -20855 772 -20838
rect 921 -20997 938 -20980
rect 672 -20997 689 -20980
rect 506 -20997 523 -20980
rect 174 -20997 191 -20980
rect 755 -20997 772 -20980
rect 921 -21139 938 -21122
rect 423 -21139 440 -21122
rect 174 -21139 191 -21122
rect 755 -21139 772 -21122
rect 921 -21281 938 -21264
rect 423 -21281 440 -21264
rect 672 -21281 689 -21264
rect 174 -21281 191 -21264
rect 755 -21281 772 -21264
rect 921 -21423 938 -21406
rect 423 -21423 440 -21406
rect 506 -21423 523 -21406
rect 174 -21423 191 -21406
rect 755 -21423 772 -21406
rect 921 -21565 938 -21548
rect 672 -21565 689 -21548
rect 506 -21565 523 -21548
rect 423 -21565 440 -21548
rect 174 -21565 191 -21548
rect 755 -21565 772 -21548
rect 921 -21707 938 -21690
rect 257 -21707 274 -21690
rect 174 -21707 191 -21690
rect 755 -21707 772 -21690
rect 921 -21849 938 -21832
rect 672 -21849 689 -21832
rect 257 -21849 274 -21832
rect 174 -21849 191 -21832
rect 755 -21849 772 -21832
rect 921 -21991 938 -21974
rect 506 -21991 523 -21974
rect 257 -21991 274 -21974
rect 174 -21991 191 -21974
rect 755 -21991 772 -21974
rect 921 -22133 938 -22116
rect 672 -22133 689 -22116
rect 506 -22133 523 -22116
rect 257 -22133 274 -22116
rect 174 -22133 191 -22116
rect 755 -22133 772 -22116
rect 921 -22275 938 -22258
rect 423 -22275 440 -22258
rect 257 -22275 274 -22258
rect 174 -22275 191 -22258
rect 755 -22275 772 -22258
rect 921 -22417 938 -22400
rect 423 -22417 440 -22400
rect 672 -22417 689 -22400
rect 257 -22417 274 -22400
rect 174 -22417 191 -22400
rect 755 -22417 772 -22400
rect 921 -22559 938 -22542
rect 423 -22559 440 -22542
rect 506 -22559 523 -22542
rect 257 -22559 274 -22542
rect 174 -22559 191 -22542
rect 755 -22559 772 -22542
rect 921 -22701 938 -22684
rect 672 -22701 689 -22684
rect 506 -22701 523 -22684
rect 423 -22701 440 -22684
rect 257 -22701 274 -22684
rect 174 -22701 191 -22684
rect 755 -22701 772 -22684
rect 921 -22843 938 -22826
rect 8 -22843 25 -22826
rect 755 -22843 772 -22826
rect 921 -22985 938 -22968
rect 8 -22985 25 -22968
rect 672 -22985 689 -22968
rect 755 -22985 772 -22968
rect 921 -23127 938 -23110
rect 8 -23127 25 -23110
rect 506 -23127 523 -23110
rect 755 -23127 772 -23110
rect 921 -23269 938 -23252
rect 8 -23269 25 -23252
rect 672 -23269 689 -23252
rect 506 -23269 523 -23252
rect 755 -23269 772 -23252
rect 921 -23411 938 -23394
rect 8 -23411 25 -23394
rect 423 -23411 440 -23394
rect 755 -23411 772 -23394
rect 921 -23553 938 -23536
rect 8 -23553 25 -23536
rect 423 -23553 440 -23536
rect 672 -23553 689 -23536
rect 755 -23553 772 -23536
rect 921 -23695 938 -23678
rect 8 -23695 25 -23678
rect 423 -23695 440 -23678
rect 506 -23695 523 -23678
rect 755 -23695 772 -23678
rect 921 -23837 938 -23820
rect 8 -23837 25 -23820
rect 672 -23837 689 -23820
rect 506 -23837 523 -23820
rect 423 -23837 440 -23820
rect 755 -23837 772 -23820
rect 921 -23979 938 -23962
rect 8 -23979 25 -23962
rect 257 -23979 274 -23962
rect 755 -23979 772 -23962
rect 921 -24121 938 -24104
rect 8 -24121 25 -24104
rect 672 -24121 689 -24104
rect 257 -24121 274 -24104
rect 755 -24121 772 -24104
rect 921 -24263 938 -24246
rect 8 -24263 25 -24246
rect 506 -24263 523 -24246
rect 257 -24263 274 -24246
rect 755 -24263 772 -24246
rect 921 -24405 938 -24388
rect 8 -24405 25 -24388
rect 672 -24405 689 -24388
rect 506 -24405 523 -24388
rect 257 -24405 274 -24388
rect 755 -24405 772 -24388
rect 921 -24547 938 -24530
rect 8 -24547 25 -24530
rect 423 -24547 440 -24530
rect 257 -24547 274 -24530
rect 755 -24547 772 -24530
rect 921 -24689 938 -24672
rect 8 -24689 25 -24672
rect 423 -24689 440 -24672
rect 672 -24689 689 -24672
rect 257 -24689 274 -24672
rect 755 -24689 772 -24672
rect 921 -24831 938 -24814
rect 8 -24831 25 -24814
rect 423 -24831 440 -24814
rect 506 -24831 523 -24814
rect 257 -24831 274 -24814
rect 755 -24831 772 -24814
rect 921 -24973 938 -24956
rect 8 -24973 25 -24956
rect 672 -24973 689 -24956
rect 506 -24973 523 -24956
rect 423 -24973 440 -24956
rect 257 -24973 274 -24956
rect 755 -24973 772 -24956
rect 921 -25115 938 -25098
rect 8 -25115 25 -25098
rect 174 -25115 191 -25098
rect 755 -25115 772 -25098
rect 921 -25257 938 -25240
rect 8 -25257 25 -25240
rect 672 -25257 689 -25240
rect 174 -25257 191 -25240
rect 755 -25257 772 -25240
rect 921 -25399 938 -25382
rect 8 -25399 25 -25382
rect 506 -25399 523 -25382
rect 174 -25399 191 -25382
rect 755 -25399 772 -25382
rect 921 -25541 938 -25524
rect 8 -25541 25 -25524
rect 672 -25541 689 -25524
rect 506 -25541 523 -25524
rect 174 -25541 191 -25524
rect 755 -25541 772 -25524
rect 921 -25683 938 -25666
rect 8 -25683 25 -25666
rect 423 -25683 440 -25666
rect 174 -25683 191 -25666
rect 755 -25683 772 -25666
rect 921 -25825 938 -25808
rect 8 -25825 25 -25808
rect 423 -25825 440 -25808
rect 672 -25825 689 -25808
rect 174 -25825 191 -25808
rect 755 -25825 772 -25808
rect 921 -25967 938 -25950
rect 8 -25967 25 -25950
rect 423 -25967 440 -25950
rect 506 -25967 523 -25950
rect 174 -25967 191 -25950
rect 755 -25967 772 -25950
rect 921 -26109 938 -26092
rect 8 -26109 25 -26092
rect 672 -26109 689 -26092
rect 506 -26109 523 -26092
rect 423 -26109 440 -26092
rect 174 -26109 191 -26092
rect 755 -26109 772 -26092
rect 921 -26251 938 -26234
rect 8 -26251 25 -26234
rect 257 -26251 274 -26234
rect 174 -26251 191 -26234
rect 755 -26251 772 -26234
rect 921 -26393 938 -26376
rect 8 -26393 25 -26376
rect 672 -26393 689 -26376
rect 257 -26393 274 -26376
rect 174 -26393 191 -26376
rect 755 -26393 772 -26376
rect 921 -26535 938 -26518
rect 8 -26535 25 -26518
rect 506 -26535 523 -26518
rect 257 -26535 274 -26518
rect 174 -26535 191 -26518
rect 755 -26535 772 -26518
rect 921 -26677 938 -26660
rect 8 -26677 25 -26660
rect 672 -26677 689 -26660
rect 506 -26677 523 -26660
rect 257 -26677 274 -26660
rect 174 -26677 191 -26660
rect 755 -26677 772 -26660
rect 921 -26819 938 -26802
rect 8 -26819 25 -26802
rect 423 -26819 440 -26802
rect 257 -26819 274 -26802
rect 174 -26819 191 -26802
rect 755 -26819 772 -26802
rect 921 -26961 938 -26944
rect 8 -26961 25 -26944
rect 423 -26961 440 -26944
rect 672 -26961 689 -26944
rect 257 -26961 274 -26944
rect 174 -26961 191 -26944
rect 755 -26961 772 -26944
rect 921 -27103 938 -27086
rect 8 -27103 25 -27086
rect 423 -27103 440 -27086
rect 506 -27103 523 -27086
rect 257 -27103 274 -27086
rect 174 -27103 191 -27086
rect 755 -27103 772 -27086
rect 921 -27245 938 -27228
rect 8 -27245 25 -27228
rect 672 -27245 689 -27228
rect 506 -27245 523 -27228
rect 423 -27245 440 -27228
rect 257 -27245 274 -27228
rect 174 -27245 191 -27228
rect 755 -27245 772 -27228
rect 921 -27387 938 -27370
rect 8 -27387 25 -27370
rect 672 -27387 689 -27370
rect 506 -27387 523 -27370
rect 423 -27387 440 -27370
rect 257 -27387 274 -27370
rect 174 -27387 191 -27370
rect 755 -27387 772 -27370
rect 921 -27529 938 -27512
rect 8 -27529 25 -27512
rect 423 -27529 440 -27512
rect 506 -27529 523 -27512
rect 257 -27529 274 -27512
rect 174 -27529 191 -27512
rect 755 -27529 772 -27512
rect 672 -27529 689 -27512
rect 921 -27671 938 -27654
rect 8 -27671 25 -27654
rect 423 -27671 440 -27654
rect 672 -27671 689 -27654
rect 257 -27671 274 -27654
rect 174 -27671 191 -27654
rect 755 -27671 772 -27654
rect 921 -27813 938 -27796
rect 8 -27813 25 -27796
rect 423 -27813 440 -27796
rect 672 -27813 689 -27796
rect 257 -27813 274 -27796
rect 174 -27813 191 -27796
rect 755 -27813 772 -27796
rect 506 -27813 523 -27796
rect 921 -27955 938 -27938
rect 8 -27955 25 -27938
rect 672 -27955 689 -27938
rect 506 -27955 523 -27938
rect 257 -27955 274 -27938
rect 174 -27955 191 -27938
rect 755 -27955 772 -27938
rect 921 -28097 938 -28080
rect 8 -28097 25 -28080
rect 506 -28097 523 -28080
rect 672 -28097 689 -28080
rect 257 -28097 274 -28080
rect 174 -28097 191 -28080
rect 755 -28097 772 -28080
rect 921 -28239 938 -28222
rect 8 -28239 25 -28222
rect 672 -28239 689 -28222
rect 257 -28239 274 -28222
rect 174 -28239 191 -28222
rect 755 -28239 772 -28222
rect 921 -28381 938 -28364
rect 8 -28381 25 -28364
rect 672 -28381 689 -28364
rect 506 -28381 523 -28364
rect 257 -28381 274 -28364
rect 174 -28381 191 -28364
rect 755 -28381 772 -28364
rect 423 -28381 440 -28364
rect 921 -28523 938 -28506
rect 8 -28523 25 -28506
rect 672 -28523 689 -28506
rect 506 -28523 523 -28506
rect 423 -28523 440 -28506
rect 174 -28523 191 -28506
rect 755 -28523 772 -28506
rect 921 -28665 938 -28648
rect 8 -28665 25 -28648
rect 423 -28665 440 -28648
rect 506 -28665 523 -28648
rect 672 -28665 689 -28648
rect 174 -28665 191 -28648
rect 755 -28665 772 -28648
rect 921 -28807 938 -28790
rect 8 -28807 25 -28790
rect 423 -28807 440 -28790
rect 672 -28807 689 -28790
rect 174 -28807 191 -28790
rect 755 -28807 772 -28790
rect 921 -28949 938 -28932
rect 8 -28949 25 -28932
rect 423 -28949 440 -28932
rect 672 -28949 689 -28932
rect 506 -28949 523 -28932
rect 174 -28949 191 -28932
rect 755 -28949 772 -28932
rect 921 -29091 938 -29074
rect 8 -29091 25 -29074
rect 672 -29091 689 -29074
rect 506 -29091 523 -29074
rect 174 -29091 191 -29074
rect 755 -29091 772 -29074
rect 921 -29233 938 -29216
rect 8 -29233 25 -29216
rect 506 -29233 523 -29216
rect 672 -29233 689 -29216
rect 174 -29233 191 -29216
rect 755 -29233 772 -29216
rect 921 -29375 938 -29358
rect 8 -29375 25 -29358
rect 672 -29375 689 -29358
rect 174 -29375 191 -29358
rect 755 -29375 772 -29358
rect 921 -29517 938 -29500
rect 257 -29517 274 -29500
rect 8 -29517 25 -29500
rect 672 -29517 689 -29500
rect 506 -29517 523 -29500
rect 423 -29517 440 -29500
rect 174 -29517 191 -29500
rect 755 -29517 772 -29500
rect 921 -29659 938 -29642
rect 8 -29659 25 -29642
rect 672 -29659 689 -29642
rect 506 -29659 523 -29642
rect 423 -29659 440 -29642
rect 257 -29659 274 -29642
rect 755 -29659 772 -29642
rect 921 -29801 938 -29784
rect 8 -29801 25 -29784
rect 423 -29801 440 -29784
rect 506 -29801 523 -29784
rect 672 -29801 689 -29784
rect 257 -29801 274 -29784
rect 755 -29801 772 -29784
rect 921 -29943 938 -29926
rect 8 -29943 25 -29926
rect 423 -29943 440 -29926
rect 672 -29943 689 -29926
rect 257 -29943 274 -29926
rect 755 -29943 772 -29926
rect 921 -30085 938 -30068
rect 8 -30085 25 -30068
rect 423 -30085 440 -30068
rect 672 -30085 689 -30068
rect 257 -30085 274 -30068
rect 506 -30085 523 -30068
rect 755 -30085 772 -30068
rect 921 -30227 938 -30210
rect 8 -30227 25 -30210
rect 672 -30227 689 -30210
rect 506 -30227 523 -30210
rect 257 -30227 274 -30210
rect 755 -30227 772 -30210
rect 921 -30369 938 -30352
rect 8 -30369 25 -30352
rect 672 -30369 689 -30352
rect 506 -30369 523 -30352
rect 257 -30369 274 -30352
rect 755 -30369 772 -30352
rect 921 -30511 938 -30494
rect 8 -30511 25 -30494
rect 672 -30511 689 -30494
rect 257 -30511 274 -30494
rect 755 -30511 772 -30494
rect 921 -30653 938 -30636
rect 8 -30653 25 -30636
rect 672 -30653 689 -30636
rect 506 -30653 523 -30636
rect 423 -30653 440 -30636
rect 257 -30653 274 -30636
rect 755 -30653 772 -30636
rect 921 -30795 938 -30778
rect 8 -30795 25 -30778
rect 672 -30795 689 -30778
rect 506 -30795 523 -30778
rect 423 -30795 440 -30778
rect 755 -30795 772 -30778
rect 921 -30937 938 -30920
rect 8 -30937 25 -30920
rect 423 -30937 440 -30920
rect 506 -30937 523 -30920
rect 672 -30937 689 -30920
rect 755 -30937 772 -30920
rect 921 -31079 938 -31062
rect 8 -31079 25 -31062
rect 423 -31079 440 -31062
rect 672 -31079 689 -31062
rect 755 -31079 772 -31062
rect 921 -31221 938 -31204
rect 8 -31221 25 -31204
rect 423 -31221 440 -31204
rect 672 -31221 689 -31204
rect 506 -31221 523 -31204
rect 755 -31221 772 -31204
rect 921 -31363 938 -31346
rect 8 -31363 25 -31346
rect 672 -31363 689 -31346
rect 506 -31363 523 -31346
rect 755 -31363 772 -31346
rect 921 -31505 938 -31488
rect 8 -31505 25 -31488
rect 672 -31505 689 -31488
rect 506 -31505 523 -31488
rect 755 -31505 772 -31488
rect 921 -31647 938 -31630
rect 8 -31647 25 -31630
rect 672 -31647 689 -31630
rect 755 -31647 772 -31630
rect 921 -31789 938 -31772
rect 8 -31789 25 -31772
rect 672 -31789 689 -31772
rect 506 -31789 523 -31772
rect 423 -31789 440 -31772
rect 257 -31789 274 -31772
rect 174 -31789 191 -31772
rect 755 -31789 772 -31772
rect 921 -31931 938 -31914
rect 672 -31931 689 -31914
rect 506 -31931 523 -31914
rect 423 -31931 440 -31914
rect 257 -31931 274 -31914
rect 174 -31931 191 -31914
rect 755 -31931 772 -31914
rect 921 -32073 938 -32056
rect 423 -32073 440 -32056
rect 506 -32073 523 -32056
rect 257 -32073 274 -32056
rect 174 -32073 191 -32056
rect 755 -32073 772 -32056
rect 672 -32073 689 -32056
rect 921 -32215 938 -32198
rect 423 -32215 440 -32198
rect 672 -32215 689 -32198
rect 257 -32215 274 -32198
rect 174 -32215 191 -32198
rect 755 -32215 772 -32198
rect 921 -32357 938 -32340
rect 423 -32357 440 -32340
rect 672 -32357 689 -32340
rect 257 -32357 274 -32340
rect 174 -32357 191 -32340
rect 755 -32357 772 -32340
rect 506 -32357 523 -32340
rect 921 -32499 938 -32482
rect 672 -32499 689 -32482
rect 506 -32499 523 -32482
rect 257 -32499 274 -32482
rect 174 -32499 191 -32482
rect 755 -32499 772 -32482
rect 921 -32641 938 -32624
rect 506 -32641 523 -32624
rect 672 -32641 689 -32624
rect 257 -32641 274 -32624
rect 174 -32641 191 -32624
rect 755 -32641 772 -32624
rect 921 -32783 938 -32766
rect 672 -32783 689 -32766
rect 257 -32783 274 -32766
rect 174 -32783 191 -32766
rect 755 -32783 772 -32766
rect 921 -32925 938 -32908
rect 672 -32925 689 -32908
rect 506 -32925 523 -32908
rect 257 -32925 274 -32908
rect 174 -32925 191 -32908
rect 755 -32925 772 -32908
rect 423 -32925 440 -32908
rect 921 -33067 938 -33050
rect 672 -33067 689 -33050
rect 506 -33067 523 -33050
rect 423 -33067 440 -33050
rect 174 -33067 191 -33050
rect 755 -33067 772 -33050
rect 921 -33209 938 -33192
rect 423 -33209 440 -33192
rect 506 -33209 523 -33192
rect 672 -33209 689 -33192
rect 174 -33209 191 -33192
rect 755 -33209 772 -33192
rect 921 -33351 938 -33334
rect 423 -33351 440 -33334
rect 672 -33351 689 -33334
rect 174 -33351 191 -33334
rect 755 -33351 772 -33334
rect 921 -33493 938 -33476
rect 423 -33493 440 -33476
rect 672 -33493 689 -33476
rect 506 -33493 523 -33476
rect 174 -33493 191 -33476
rect 755 -33493 772 -33476
rect 921 -33635 938 -33618
rect 672 -33635 689 -33618
rect 506 -33635 523 -33618
rect 174 -33635 191 -33618
rect 755 -33635 772 -33618
rect 921 -33777 938 -33760
rect 506 -33777 523 -33760
rect 672 -33777 689 -33760
rect 174 -33777 191 -33760
rect 755 -33777 772 -33760
rect 921 -33919 938 -33902
rect 672 -33919 689 -33902
rect 174 -33919 191 -33902
rect 755 -33919 772 -33902
rect 921 -34061 938 -34044
rect 257 -34061 274 -34044
rect 672 -34061 689 -34044
rect 506 -34061 523 -34044
rect 423 -34061 440 -34044
rect 174 -34061 191 -34044
rect 755 -34061 772 -34044
rect 921 -34203 938 -34186
rect 672 -34203 689 -34186
rect 506 -34203 523 -34186
rect 423 -34203 440 -34186
rect 257 -34203 274 -34186
rect 755 -34203 772 -34186
rect 921 -34345 938 -34328
rect 423 -34345 440 -34328
rect 506 -34345 523 -34328
rect 672 -34345 689 -34328
rect 257 -34345 274 -34328
rect 755 -34345 772 -34328
rect 921 -34487 938 -34470
rect 423 -34487 440 -34470
rect 672 -34487 689 -34470
rect 257 -34487 274 -34470
rect 755 -34487 772 -34470
rect 921 -34629 938 -34612
rect 423 -34629 440 -34612
rect 672 -34629 689 -34612
rect 257 -34629 274 -34612
rect 506 -34629 523 -34612
rect 755 -34629 772 -34612
rect 921 -34771 938 -34754
rect 672 -34771 689 -34754
rect 506 -34771 523 -34754
rect 257 -34771 274 -34754
rect 755 -34771 772 -34754
rect 921 -34913 938 -34896
rect 672 -34913 689 -34896
rect 506 -34913 523 -34896
rect 257 -34913 274 -34896
rect 755 -34913 772 -34896
rect 921 -35055 938 -35038
rect 672 -35055 689 -35038
rect 257 -35055 274 -35038
rect 755 -35055 772 -35038
rect 921 -35197 938 -35180
rect 672 -35197 689 -35180
rect 506 -35197 523 -35180
rect 423 -35197 440 -35180
rect 257 -35197 274 -35180
rect 755 -35197 772 -35180
rect 921 -35339 938 -35322
rect 672 -35339 689 -35322
rect 506 -35339 523 -35322
rect 423 -35339 440 -35322
rect 755 -35339 772 -35322
rect 921 -35481 938 -35464
rect 423 -35481 440 -35464
rect 506 -35481 523 -35464
rect 672 -35481 689 -35464
rect 755 -35481 772 -35464
rect 921 -35623 938 -35606
rect 423 -35623 440 -35606
rect 672 -35623 689 -35606
rect 755 -35623 772 -35606
rect 921 -35765 938 -35748
rect 423 -35765 440 -35748
rect 672 -35765 689 -35748
rect 506 -35765 523 -35748
rect 755 -35765 772 -35748
rect 921 -35907 938 -35890
rect 672 -35907 689 -35890
rect 506 -35907 523 -35890
rect 755 -35907 772 -35890
rect 921 -36049 938 -36032
rect 672 -36049 689 -36032
rect 506 -36049 523 -36032
rect 755 -36049 772 -36032
rect 921 -36191 938 -36174
rect 672 -36191 689 -36174
rect 755 -36191 772 -36174
rect 921 -36333 938 -36316
rect 921 -36475 938 -36458
rect 921 -36617 938 -36600
rect 755 -36617 772 -36600
rect 921 -36759 938 -36742
rect 672 -36759 689 -36742
rect 921 -36901 938 -36884
rect 672 -36901 689 -36884
rect 755 -36901 772 -36884
rect 921 -37043 938 -37026
rect 506 -37043 523 -37026
rect 921 -37185 938 -37168
rect 506 -37185 523 -37168
rect 755 -37185 772 -37168
rect 921 -37327 938 -37310
rect 672 -37327 689 -37310
rect 506 -37327 523 -37310
rect 921 -37469 938 -37452
rect 672 -37469 689 -37452
rect 506 -37469 523 -37452
rect 755 -37469 772 -37452
rect 921 -37611 938 -37594
rect 423 -37611 440 -37594
rect 921 -37753 938 -37736
rect 423 -37753 440 -37736
rect 755 -37753 772 -37736
rect 921 -37895 938 -37878
rect 423 -37895 440 -37878
rect 672 -37895 689 -37878
rect 921 -38037 938 -38020
rect 672 -38037 689 -38020
rect 423 -38037 440 -38020
rect 755 -38037 772 -38020
rect 921 -38179 938 -38162
rect 423 -38179 440 -38162
rect 506 -38179 523 -38162
rect 921 -38321 938 -38304
rect 423 -38321 440 -38304
rect 506 -38321 523 -38304
rect 755 -38321 772 -38304
rect 921 -38463 938 -38446
rect 423 -38463 440 -38446
rect 672 -38463 689 -38446
rect 506 -38463 523 -38446
rect 921 -38605 938 -38588
rect 672 -38605 689 -38588
rect 506 -38605 523 -38588
rect 423 -38605 440 -38588
rect 755 -38605 772 -38588
rect 257 -38747 274 -38730
rect 921 -38747 938 -38730
rect 921 -38889 938 -38872
rect 257 -38889 274 -38872
rect 755 -38889 772 -38872
rect 921 -39031 938 -39014
rect 672 -39031 689 -39014
rect 257 -39031 274 -39014
rect 921 -39173 938 -39156
rect 672 -39173 689 -39156
rect 257 -39173 274 -39156
rect 755 -39173 772 -39156
rect 921 -39315 938 -39298
rect 506 -39315 523 -39298
rect 257 -39315 274 -39298
rect 921 -39457 938 -39440
rect 506 -39457 523 -39440
rect 257 -39457 274 -39440
rect 755 -39457 772 -39440
rect 921 -39599 938 -39582
rect 672 -39599 689 -39582
rect 506 -39599 523 -39582
rect 257 -39599 274 -39582
rect 921 -39741 938 -39724
rect 672 -39741 689 -39724
rect 506 -39741 523 -39724
rect 257 -39741 274 -39724
rect 755 -39741 772 -39724
rect 921 -39883 938 -39866
rect 423 -39883 440 -39866
rect 257 -39883 274 -39866
rect 921 -40025 938 -40008
rect 423 -40025 440 -40008
rect 257 -40025 274 -40008
rect 755 -40025 772 -40008
rect 921 -40167 938 -40150
rect 423 -40167 440 -40150
rect 672 -40167 689 -40150
rect 257 -40167 274 -40150
rect 921 -40309 938 -40292
rect 672 -40309 689 -40292
rect 423 -40309 440 -40292
rect 257 -40309 274 -40292
rect 755 -40309 772 -40292
rect 921 -40451 938 -40434
rect 423 -40451 440 -40434
rect 506 -40451 523 -40434
rect 257 -40451 274 -40434
rect 921 -40593 938 -40576
rect 423 -40593 440 -40576
rect 506 -40593 523 -40576
rect 257 -40593 274 -40576
rect 755 -40593 772 -40576
rect 921 -40735 938 -40718
rect 423 -40735 440 -40718
rect 672 -40735 689 -40718
rect 506 -40735 523 -40718
rect 257 -40735 274 -40718
rect 921 -40877 938 -40860
rect 672 -40877 689 -40860
rect 506 -40877 523 -40860
rect 423 -40877 440 -40860
rect 257 -40877 274 -40860
rect 755 -40877 772 -40860
rect 174 -41019 191 -41002
rect 921 -41019 938 -41002
rect 921 -41161 938 -41144
rect 174 -41161 191 -41144
rect 755 -41161 772 -41144
rect 921 -41303 938 -41286
rect 672 -41303 689 -41286
rect 174 -41303 191 -41286
rect 921 -41445 938 -41428
rect 672 -41445 689 -41428
rect 174 -41445 191 -41428
rect 755 -41445 772 -41428
rect 921 -41587 938 -41570
rect 506 -41587 523 -41570
rect 174 -41587 191 -41570
rect 921 -41729 938 -41712
rect 506 -41729 523 -41712
rect 174 -41729 191 -41712
rect 755 -41729 772 -41712
rect 921 -41871 938 -41854
rect 672 -41871 689 -41854
rect 506 -41871 523 -41854
rect 174 -41871 191 -41854
rect 921 -42013 938 -41996
rect 672 -42013 689 -41996
rect 506 -42013 523 -41996
rect 174 -42013 191 -41996
rect 755 -42013 772 -41996
rect 921 -42155 938 -42138
rect 423 -42155 440 -42138
rect 174 -42155 191 -42138
rect 921 -42297 938 -42280
rect 423 -42297 440 -42280
rect 174 -42297 191 -42280
rect 755 -42297 772 -42280
rect 921 -42439 938 -42422
rect 423 -42439 440 -42422
rect 672 -42439 689 -42422
rect 174 -42439 191 -42422
rect 921 -42581 938 -42564
rect 672 -42581 689 -42564
rect 423 -42581 440 -42564
rect 174 -42581 191 -42564
rect 755 -42581 772 -42564
rect 921 -42723 938 -42706
rect 423 -42723 440 -42706
rect 506 -42723 523 -42706
rect 174 -42723 191 -42706
rect 921 -42865 938 -42848
rect 423 -42865 440 -42848
rect 506 -42865 523 -42848
rect 174 -42865 191 -42848
rect 755 -42865 772 -42848
rect 921 -43007 938 -42990
rect 423 -43007 440 -42990
rect 672 -43007 689 -42990
rect 506 -43007 523 -42990
rect 174 -43007 191 -42990
rect 921 -43149 938 -43132
rect 672 -43149 689 -43132
rect 506 -43149 523 -43132
rect 423 -43149 440 -43132
rect 174 -43149 191 -43132
rect 755 -43149 772 -43132
rect 921 -43291 938 -43274
rect 257 -43291 274 -43274
rect 174 -43291 191 -43274
rect 921 -43433 938 -43416
rect 257 -43433 274 -43416
rect 174 -43433 191 -43416
rect 755 -43433 772 -43416
rect 921 -43575 938 -43558
rect 672 -43575 689 -43558
rect 257 -43575 274 -43558
rect 174 -43575 191 -43558
rect 921 -43717 938 -43700
rect 672 -43717 689 -43700
rect 257 -43717 274 -43700
rect 174 -43717 191 -43700
rect 755 -43717 772 -43700
rect 921 -43859 938 -43842
rect 506 -43859 523 -43842
rect 257 -43859 274 -43842
rect 174 -43859 191 -43842
rect 921 -44001 938 -43984
rect 506 -44001 523 -43984
rect 257 -44001 274 -43984
rect 174 -44001 191 -43984
rect 755 -44001 772 -43984
rect 921 -44143 938 -44126
rect 672 -44143 689 -44126
rect 506 -44143 523 -44126
rect 257 -44143 274 -44126
rect 174 -44143 191 -44126
rect 921 -44285 938 -44268
rect 672 -44285 689 -44268
rect 506 -44285 523 -44268
rect 257 -44285 274 -44268
rect 174 -44285 191 -44268
rect 755 -44285 772 -44268
rect 921 -44427 938 -44410
rect 423 -44427 440 -44410
rect 257 -44427 274 -44410
rect 174 -44427 191 -44410
rect 921 -44569 938 -44552
rect 423 -44569 440 -44552
rect 257 -44569 274 -44552
rect 174 -44569 191 -44552
rect 755 -44569 772 -44552
rect 921 -44711 938 -44694
rect 423 -44711 440 -44694
rect 672 -44711 689 -44694
rect 257 -44711 274 -44694
rect 174 -44711 191 -44694
rect 921 -44853 938 -44836
rect 672 -44853 689 -44836
rect 423 -44853 440 -44836
rect 257 -44853 274 -44836
rect 174 -44853 191 -44836
rect 755 -44853 772 -44836
rect 921 -44995 938 -44978
rect 423 -44995 440 -44978
rect 506 -44995 523 -44978
rect 257 -44995 274 -44978
rect 174 -44995 191 -44978
rect 921 -45137 938 -45120
rect 423 -45137 440 -45120
rect 506 -45137 523 -45120
rect 257 -45137 274 -45120
rect 174 -45137 191 -45120
rect 755 -45137 772 -45120
rect 921 -45279 938 -45262
rect 423 -45279 440 -45262
rect 672 -45279 689 -45262
rect 506 -45279 523 -45262
rect 257 -45279 274 -45262
rect 174 -45279 191 -45262
rect 921 -45421 938 -45404
rect 672 -45421 689 -45404
rect 506 -45421 523 -45404
rect 423 -45421 440 -45404
rect 257 -45421 274 -45404
rect 174 -45421 191 -45404
rect 755 -45421 772 -45404
rect 8 -45563 25 -45546
rect 921 -45563 938 -45546
rect 921 -45705 938 -45688
rect 8 -45705 25 -45688
rect 755 -45705 772 -45688
rect 921 -45847 938 -45830
rect 8 -45847 25 -45830
rect 672 -45847 689 -45830
rect 921 -45989 938 -45972
rect 8 -45989 25 -45972
rect 672 -45989 689 -45972
rect 755 -45989 772 -45972
rect 921 -46131 938 -46114
rect 8 -46131 25 -46114
rect 506 -46131 523 -46114
rect 921 -46273 938 -46256
rect 8 -46273 25 -46256
rect 506 -46273 523 -46256
rect 755 -46273 772 -46256
rect 921 -46415 938 -46398
rect 8 -46415 25 -46398
rect 672 -46415 689 -46398
rect 506 -46415 523 -46398
rect 921 -46557 938 -46540
rect 8 -46557 25 -46540
rect 672 -46557 689 -46540
rect 506 -46557 523 -46540
rect 755 -46557 772 -46540
rect 921 -46699 938 -46682
rect 8 -46699 25 -46682
rect 423 -46699 440 -46682
rect 921 -46841 938 -46824
rect 8 -46841 25 -46824
rect 423 -46841 440 -46824
rect 755 -46841 772 -46824
rect 921 -46983 938 -46966
rect 8 -46983 25 -46966
rect 423 -46983 440 -46966
rect 672 -46983 689 -46966
rect 921 -47125 938 -47108
rect 8 -47125 25 -47108
rect 672 -47125 689 -47108
rect 423 -47125 440 -47108
rect 755 -47125 772 -47108
rect 921 -47267 938 -47250
rect 8 -47267 25 -47250
rect 423 -47267 440 -47250
rect 506 -47267 523 -47250
rect 921 -47409 938 -47392
rect 8 -47409 25 -47392
rect 423 -47409 440 -47392
rect 506 -47409 523 -47392
rect 755 -47409 772 -47392
rect 921 -47551 938 -47534
rect 8 -47551 25 -47534
rect 423 -47551 440 -47534
rect 672 -47551 689 -47534
rect 506 -47551 523 -47534
rect 921 -47693 938 -47676
rect 8 -47693 25 -47676
rect 672 -47693 689 -47676
rect 506 -47693 523 -47676
rect 423 -47693 440 -47676
rect 755 -47693 772 -47676
rect 921 -47835 938 -47818
rect 8 -47835 25 -47818
rect 257 -47835 274 -47818
rect 921 -47977 938 -47960
rect 8 -47977 25 -47960
rect 257 -47977 274 -47960
rect 755 -47977 772 -47960
rect 921 -48119 938 -48102
rect 8 -48119 25 -48102
rect 672 -48119 689 -48102
rect 257 -48119 274 -48102
rect 921 -48261 938 -48244
rect 8 -48261 25 -48244
rect 672 -48261 689 -48244
rect 257 -48261 274 -48244
rect 755 -48261 772 -48244
rect 921 -48403 938 -48386
rect 8 -48403 25 -48386
rect 506 -48403 523 -48386
rect 257 -48403 274 -48386
rect 921 -48545 938 -48528
rect 8 -48545 25 -48528
rect 506 -48545 523 -48528
rect 257 -48545 274 -48528
rect 755 -48545 772 -48528
rect 921 -48687 938 -48670
rect 8 -48687 25 -48670
rect 672 -48687 689 -48670
rect 506 -48687 523 -48670
rect 257 -48687 274 -48670
rect 921 -48829 938 -48812
rect 8 -48829 25 -48812
rect 672 -48829 689 -48812
rect 506 -48829 523 -48812
rect 257 -48829 274 -48812
rect 755 -48829 772 -48812
rect 921 -48971 938 -48954
rect 8 -48971 25 -48954
rect 423 -48971 440 -48954
rect 257 -48971 274 -48954
rect 921 -49113 938 -49096
rect 8 -49113 25 -49096
rect 423 -49113 440 -49096
rect 257 -49113 274 -49096
rect 755 -49113 772 -49096
rect 921 -49255 938 -49238
rect 8 -49255 25 -49238
rect 423 -49255 440 -49238
rect 672 -49255 689 -49238
rect 257 -49255 274 -49238
rect 921 -49397 938 -49380
rect 8 -49397 25 -49380
rect 672 -49397 689 -49380
rect 423 -49397 440 -49380
rect 257 -49397 274 -49380
rect 755 -49397 772 -49380
rect 921 -49539 938 -49522
rect 8 -49539 25 -49522
rect 423 -49539 440 -49522
rect 506 -49539 523 -49522
rect 257 -49539 274 -49522
rect 921 -49681 938 -49664
rect 8 -49681 25 -49664
rect 423 -49681 440 -49664
rect 506 -49681 523 -49664
rect 257 -49681 274 -49664
rect 755 -49681 772 -49664
rect 921 -49823 938 -49806
rect 8 -49823 25 -49806
rect 423 -49823 440 -49806
rect 672 -49823 689 -49806
rect 506 -49823 523 -49806
rect 257 -49823 274 -49806
rect 921 -49965 938 -49948
rect 8 -49965 25 -49948
rect 672 -49965 689 -49948
rect 506 -49965 523 -49948
rect 423 -49965 440 -49948
rect 257 -49965 274 -49948
rect 755 -49965 772 -49948
rect 921 -50107 938 -50090
rect 8 -50107 25 -50090
rect 174 -50107 191 -50090
rect 921 -50249 938 -50232
rect 8 -50249 25 -50232
rect 174 -50249 191 -50232
rect 755 -50249 772 -50232
rect 921 -50391 938 -50374
rect 8 -50391 25 -50374
rect 672 -50391 689 -50374
rect 174 -50391 191 -50374
rect 921 -50533 938 -50516
rect 8 -50533 25 -50516
rect 672 -50533 689 -50516
rect 174 -50533 191 -50516
rect 755 -50533 772 -50516
rect 921 -50675 938 -50658
rect 8 -50675 25 -50658
rect 506 -50675 523 -50658
rect 174 -50675 191 -50658
rect 921 -50817 938 -50800
rect 8 -50817 25 -50800
rect 506 -50817 523 -50800
rect 174 -50817 191 -50800
rect 755 -50817 772 -50800
rect 921 -50959 938 -50942
rect 8 -50959 25 -50942
rect 672 -50959 689 -50942
rect 506 -50959 523 -50942
rect 174 -50959 191 -50942
rect 921 -51101 938 -51084
rect 8 -51101 25 -51084
rect 672 -51101 689 -51084
rect 506 -51101 523 -51084
rect 174 -51101 191 -51084
rect 755 -51101 772 -51084
rect 921 -51243 938 -51226
rect 8 -51243 25 -51226
rect 423 -51243 440 -51226
rect 174 -51243 191 -51226
rect 921 -51385 938 -51368
rect 8 -51385 25 -51368
rect 423 -51385 440 -51368
rect 174 -51385 191 -51368
rect 755 -51385 772 -51368
rect 921 -51527 938 -51510
rect 8 -51527 25 -51510
rect 423 -51527 440 -51510
rect 672 -51527 689 -51510
rect 174 -51527 191 -51510
rect 921 -51669 938 -51652
rect 8 -51669 25 -51652
rect 672 -51669 689 -51652
rect 423 -51669 440 -51652
rect 174 -51669 191 -51652
rect 755 -51669 772 -51652
rect 921 -51811 938 -51794
rect 8 -51811 25 -51794
rect 423 -51811 440 -51794
rect 506 -51811 523 -51794
rect 174 -51811 191 -51794
rect 921 -51953 938 -51936
rect 8 -51953 25 -51936
rect 423 -51953 440 -51936
rect 506 -51953 523 -51936
rect 174 -51953 191 -51936
rect 755 -51953 772 -51936
rect 921 -52095 938 -52078
rect 8 -52095 25 -52078
rect 423 -52095 440 -52078
rect 672 -52095 689 -52078
rect 506 -52095 523 -52078
rect 174 -52095 191 -52078
rect 921 -52237 938 -52220
rect 8 -52237 25 -52220
rect 672 -52237 689 -52220
rect 506 -52237 523 -52220
rect 423 -52237 440 -52220
rect 174 -52237 191 -52220
rect 755 -52237 772 -52220
rect 921 -52379 938 -52362
rect 8 -52379 25 -52362
rect 257 -52379 274 -52362
rect 174 -52379 191 -52362
rect 921 -52521 938 -52504
rect 8 -52521 25 -52504
rect 257 -52521 274 -52504
rect 174 -52521 191 -52504
rect 755 -52521 772 -52504
rect 921 -52663 938 -52646
rect 8 -52663 25 -52646
rect 672 -52663 689 -52646
rect 257 -52663 274 -52646
rect 174 -52663 191 -52646
rect 921 -52805 938 -52788
rect 8 -52805 25 -52788
rect 672 -52805 689 -52788
rect 257 -52805 274 -52788
rect 174 -52805 191 -52788
rect 755 -52805 772 -52788
rect 921 -52947 938 -52930
rect 8 -52947 25 -52930
rect 506 -52947 523 -52930
rect 257 -52947 274 -52930
rect 174 -52947 191 -52930
rect 921 -53089 938 -53072
rect 8 -53089 25 -53072
rect 506 -53089 523 -53072
rect 257 -53089 274 -53072
rect 174 -53089 191 -53072
rect 755 -53089 772 -53072
rect 921 -53231 938 -53214
rect 8 -53231 25 -53214
rect 672 -53231 689 -53214
rect 506 -53231 523 -53214
rect 257 -53231 274 -53214
rect 174 -53231 191 -53214
rect 921 -53373 938 -53356
rect 8 -53373 25 -53356
rect 672 -53373 689 -53356
rect 506 -53373 523 -53356
rect 257 -53373 274 -53356
rect 174 -53373 191 -53356
rect 755 -53373 772 -53356
rect 921 -53515 938 -53498
rect 8 -53515 25 -53498
rect 423 -53515 440 -53498
rect 257 -53515 274 -53498
rect 174 -53515 191 -53498
rect 921 -53657 938 -53640
rect 8 -53657 25 -53640
rect 423 -53657 440 -53640
rect 257 -53657 274 -53640
rect 174 -53657 191 -53640
rect 755 -53657 772 -53640
rect 921 -53799 938 -53782
rect 8 -53799 25 -53782
rect 423 -53799 440 -53782
rect 672 -53799 689 -53782
rect 257 -53799 274 -53782
rect 174 -53799 191 -53782
rect 921 -53941 938 -53924
rect 8 -53941 25 -53924
rect 672 -53941 689 -53924
rect 423 -53941 440 -53924
rect 257 -53941 274 -53924
rect 174 -53941 191 -53924
rect 755 -53941 772 -53924
rect 921 -54083 938 -54066
rect 8 -54083 25 -54066
rect 423 -54083 440 -54066
rect 506 -54083 523 -54066
rect 257 -54083 274 -54066
rect 174 -54083 191 -54066
rect 921 -54225 938 -54208
rect 8 -54225 25 -54208
rect 423 -54225 440 -54208
rect 506 -54225 523 -54208
rect 257 -54225 274 -54208
rect 174 -54225 191 -54208
rect 755 -54225 772 -54208
rect 921 -54367 938 -54350
rect 8 -54367 25 -54350
rect 423 -54367 440 -54350
rect 672 -54367 689 -54350
rect 506 -54367 523 -54350
rect 257 -54367 274 -54350
rect 174 -54367 191 -54350
rect 8 -54509 25 -54492
rect 672 -54509 689 -54492
rect 506 -54509 523 -54492
rect 423 -54509 440 -54492
rect 257 -54509 274 -54492
rect 174 -54509 191 -54492
rect 755 -54509 772 -54492
rect 921 -54793 938 -54776
rect 921 -54935 938 -54918
rect 755 -55077 772 -55060
rect 921 -55219 938 -55202
rect 672 -55219 689 -55202
rect 755 -55219 772 -55202
rect 921 -55361 938 -55344
rect 672 -55361 689 -55344
rect 921 -55503 938 -55486
rect 672 -55503 689 -55486
rect 755 -55503 772 -55486
rect 921 -55645 938 -55628
rect 506 -55645 523 -55628
rect 755 -55645 772 -55628
rect 921 -55787 938 -55770
rect 672 -55787 689 -55770
rect 506 -55787 523 -55770
rect 755 -55787 772 -55770
rect 921 -55929 938 -55912
rect 672 -55929 689 -55912
rect 506 -55929 523 -55912
rect 755 -55929 772 -55912
rect 921 -56071 938 -56054
rect 423 -56071 440 -56054
rect 755 -56071 772 -56054
rect 921 -56213 938 -56196
rect 423 -56213 440 -56196
rect 672 -56213 689 -56196
rect 921 -56355 938 -56338
rect 672 -56355 689 -56338
rect 423 -56355 440 -56338
rect 506 -56355 523 -56338
rect 755 -56355 772 -56338
rect 921 -56497 938 -56480
rect 423 -56497 440 -56480
rect 506 -56497 523 -56480
rect 672 -56497 689 -56480
rect 755 -56497 772 -56480
rect 921 -56639 938 -56622
rect 672 -56639 689 -56622
rect 506 -56639 523 -56622
rect 423 -56639 440 -56622
rect 257 -56639 274 -56622
rect 755 -56639 772 -56622
rect 921 -56781 938 -56764
rect 672 -56781 689 -56764
rect 257 -56781 274 -56764
rect 755 -56781 772 -56764
rect 506 -56923 523 -56906
rect 257 -56923 274 -56906
rect 755 -56923 772 -56906
rect 921 -57065 938 -57048
rect 672 -57065 689 -57048
rect 506 -57065 523 -57048
rect 257 -57065 274 -57048
rect 755 -57065 772 -57048
rect 921 -57207 938 -57190
rect 423 -57207 440 -57190
rect 672 -57207 689 -57190
rect 257 -57207 274 -57190
rect 921 -57349 938 -57332
rect 672 -57349 689 -57332
rect 423 -57349 440 -57332
rect 257 -57349 274 -57332
rect 506 -57349 523 -57332
rect 755 -57349 772 -57332
rect 921 -57491 938 -57474
rect 423 -57491 440 -57474
rect 506 -57491 523 -57474
rect 672 -57491 689 -57474
rect 257 -57491 274 -57474
rect 755 -57491 772 -57474
rect 921 -57633 938 -57616
rect 174 -57633 191 -57616
rect 755 -57633 772 -57616
rect 921 -57775 938 -57758
rect 672 -57775 689 -57758
rect 506 -57775 523 -57758
rect 174 -57775 191 -57758
rect 755 -57775 772 -57758
rect 921 -57917 938 -57900
rect 672 -57917 689 -57900
rect 506 -57917 523 -57900
rect 174 -57917 191 -57900
rect 755 -57917 772 -57900
rect 921 -58059 938 -58042
rect 423 -58059 440 -58042
rect 672 -58059 689 -58042
rect 174 -58059 191 -58042
rect 755 -58059 772 -58042
rect 423 -58201 440 -58184
rect 506 -58201 523 -58184
rect 174 -58201 191 -58184
rect 755 -58201 772 -58184
rect 921 -58343 938 -58326
rect 672 -58343 689 -58326
rect 506 -58343 523 -58326
rect 423 -58343 440 -58326
rect 257 -58343 274 -58326
rect 174 -58343 191 -58326
rect 921 -58485 938 -58468
rect 672 -58485 689 -58468
rect 257 -58485 274 -58468
rect 174 -58485 191 -58468
rect 755 -58485 772 -58468
rect 921 -58627 938 -58610
rect 506 -58627 523 -58610
rect 672 -58627 689 -58610
rect 257 -58627 274 -58610
rect 174 -58627 191 -58610
rect 755 -58627 772 -58610
rect 921 -58769 938 -58752
rect 423 -58769 440 -58752
rect 257 -58769 274 -58752
rect 174 -58769 191 -58752
rect 755 -58769 772 -58752
rect 921 -58911 938 -58894
rect 506 -58911 523 -58894
rect 672 -58911 689 -58894
rect 423 -58911 440 -58894
rect 257 -58911 274 -58894
rect 174 -58911 191 -58894
rect 755 -58911 772 -58894
rect 8 -59053 25 -59036
rect 423 -59053 440 -59036
rect 672 -59053 689 -59036
rect 506 -59053 523 -59036
rect 257 -59053 274 -59036
rect 174 -59053 191 -59036
rect 921 -59195 938 -59178
rect 8 -59195 25 -59178
rect 672 -59195 689 -59178
rect 755 -59195 772 -59178
rect 921 -59337 938 -59320
rect 8 -59337 25 -59320
rect 672 -59337 689 -59320
rect 506 -59337 523 -59320
rect 921 -59479 938 -59462
rect 8 -59479 25 -59462
rect 672 -59479 689 -59462
rect 506 -59479 523 -59462
rect 423 -59479 440 -59462
rect 755 -59479 772 -59462
rect 921 -59621 938 -59604
rect 8 -59621 25 -59604
rect 423 -59621 440 -59604
rect 672 -59621 689 -59604
rect 506 -59621 523 -59604
rect 921 -59763 938 -59746
rect 8 -59763 25 -59746
rect 423 -59763 440 -59746
rect 506 -59763 523 -59746
rect 672 -59763 689 -59746
rect 755 -59763 772 -59746
rect 921 -59905 938 -59888
rect 8 -59905 25 -59888
rect 672 -59905 689 -59888
rect 257 -59905 274 -59888
rect 755 -59905 772 -59888
rect 921 -60047 938 -60030
rect 8 -60047 25 -60030
rect 672 -60047 689 -60030
rect 506 -60047 523 -60030
rect 257 -60047 274 -60030
rect 755 -60047 772 -60030
rect 921 -60189 938 -60172
rect 8 -60189 25 -60172
rect 672 -60189 689 -60172
rect 506 -60189 523 -60172
rect 423 -60189 440 -60172
rect 257 -60189 274 -60172
rect 921 -60331 938 -60314
rect 8 -60331 25 -60314
rect 423 -60331 440 -60314
rect 672 -60331 689 -60314
rect 257 -60331 274 -60314
rect 755 -60331 772 -60314
rect 921 -60473 938 -60456
rect 8 -60473 25 -60456
rect 423 -60473 440 -60456
rect 506 -60473 523 -60456
rect 672 -60473 689 -60456
rect 257 -60473 274 -60456
rect 921 -60615 938 -60598
rect 8 -60615 25 -60598
rect 672 -60615 689 -60598
rect 506 -60615 523 -60598
rect 423 -60615 440 -60598
rect 257 -60615 274 -60598
rect 174 -60615 191 -60598
rect 755 -60615 772 -60598
rect 8 -60757 25 -60740
rect 672 -60757 689 -60740
rect 174 -60757 191 -60740
rect 755 -60757 772 -60740
rect 921 -60899 938 -60882
rect 8 -60899 25 -60882
rect 506 -60899 523 -60882
rect 174 -60899 191 -60882
rect 755 -60899 772 -60882
rect 8 -61041 25 -61024
rect 672 -61041 689 -61024
rect 506 -61041 523 -61024
rect 423 -61041 440 -61024
rect 174 -61041 191 -61024
rect 755 -61041 772 -61024
rect 921 -61183 938 -61166
rect 8 -61183 25 -61166
rect 423 -61183 440 -61166
rect 672 -61183 689 -61166
rect 174 -61183 191 -61166
rect 755 -61183 772 -61166
rect 921 -61325 938 -61308
rect 8 -61325 25 -61308
rect 672 -61325 689 -61308
rect 423 -61325 440 -61308
rect 174 -61325 191 -61308
rect 755 -61325 772 -61308
rect 506 -61325 523 -61308
rect 8 -61467 25 -61450
rect 423 -61467 440 -61450
rect 672 -61467 689 -61450
rect 506 -61467 523 -61450
rect 174 -61467 191 -61450
rect 755 -61467 772 -61450
rect 8 -61609 25 -61592
rect 257 -61609 274 -61592
rect 174 -61609 191 -61592
rect 755 -61609 772 -61592
rect 8 -61751 25 -61734
rect 672 -61751 689 -61734
rect 257 -61751 274 -61734
rect 174 -61751 191 -61734
rect 755 -61751 772 -61734
rect 8 -61893 25 -61876
rect 506 -61893 523 -61876
rect 257 -61893 274 -61876
rect 174 -61893 191 -61876
rect 755 -61893 772 -61876
rect 921 -62035 938 -62018
rect 8 -62035 25 -62018
rect 506 -62035 523 -62018
rect 672 -62035 689 -62018
rect 257 -62035 274 -62018
rect 174 -62035 191 -62018
rect 755 -62035 772 -62018
rect 8 -62177 25 -62160
rect 672 -62177 689 -62160
rect 506 -62177 523 -62160
rect 257 -62177 274 -62160
rect 174 -62177 191 -62160
rect 755 -62177 772 -62160
rect 423 -62177 440 -62160
rect 921 -62319 938 -62302
rect 8 -62319 25 -62302
rect 423 -62319 440 -62302
rect 257 -62319 274 -62302
rect 174 -62319 191 -62302
rect 755 -62319 772 -62302
rect 921 -62461 938 -62444
rect 8 -62461 25 -62444
rect 423 -62461 440 -62444
rect 672 -62461 689 -62444
rect 257 -62461 274 -62444
rect 174 -62461 191 -62444
rect 8 -62603 25 -62586
rect 672 -62603 689 -62586
rect 423 -62603 440 -62586
rect 257 -62603 274 -62586
rect 174 -62603 191 -62586
rect 755 -62603 772 -62586
rect 506 -62603 523 -62586
rect 921 -62745 938 -62728
rect 8 -62745 25 -62728
rect 423 -62745 440 -62728
rect 506 -62745 523 -62728
rect 257 -62745 274 -62728
rect 174 -62745 191 -62728
rect 755 -62745 772 -62728
rect 921 -62887 938 -62870
rect 8 -62887 25 -62870
rect 423 -62887 440 -62870
rect 506 -62887 523 -62870
rect 257 -62887 274 -62870
rect 174 -62887 191 -62870
rect 755 -62887 772 -62870
rect 921 -63029 938 -63012
rect 8 -63029 25 -63012
rect 423 -63029 440 -63012
rect 672 -63029 689 -63012
rect 506 -63029 523 -63012
rect 257 -63029 274 -63012
rect 174 -63029 191 -63012
rect 921 -63171 938 -63154
rect 8 -63171 25 -63154
rect 672 -63171 689 -63154
rect 506 -63171 523 -63154
rect 423 -63171 440 -63154
rect 257 -63171 274 -63154
rect 174 -63171 191 -63154
rect 755 -63171 772 -63154
rect 8 -63313 25 -63296
rect 672 -63313 689 -63296
rect 506 -63313 523 -63296
rect 423 -63313 440 -63296
rect 257 -63313 274 -63296
rect 174 -63313 191 -63296
rect 755 -63313 772 -63296
rect 921 -63455 938 -63438
rect 8 -63455 25 -63438
rect 672 -63455 689 -63438
rect 506 -63455 523 -63438
rect 423 -63455 440 -63438
rect 257 -63455 274 -63438
rect 174 -63455 191 -63438
rect 755 -63455 772 -63438
rect 921 -63597 938 -63580
rect 8 -63597 25 -63580
rect 672 -63597 689 -63580
rect 506 -63597 523 -63580
rect 423 -63597 440 -63580
rect 257 -63597 274 -63580
rect 174 -63597 191 -63580
rect 755 -63597 772 -63580
rect 921 -63739 938 -63722
rect 8 -63739 25 -63722
rect 672 -63739 689 -63722
rect 506 -63739 523 -63722
rect 423 -63739 440 -63722
rect 257 -63739 274 -63722
rect 174 -63739 191 -63722
rect 755 -63739 772 -63722
rect 921 -63881 938 -63864
rect 8 -63881 25 -63864
rect 672 -63881 689 -63864
rect 506 -63881 523 -63864
rect 423 -63881 440 -63864
rect 257 -63881 274 -63864
rect 174 -63881 191 -63864
rect 755 -63881 772 -63864
rect 8 -64023 25 -64006
rect 672 -64023 689 -64006
rect 506 -64023 523 -64006
rect 423 -64023 440 -64006
rect 257 -64023 274 -64006
rect 174 -64023 191 -64006
rect 755 -64023 772 -64006
rect 921 -64165 938 -64148
rect 8 -64165 25 -64148
rect 672 -64165 689 -64148
rect 506 -64165 523 -64148
rect 423 -64165 440 -64148
rect 257 -64165 274 -64148
rect 174 -64165 191 -64148
rect 921 -64307 938 -64290
rect 8 -64307 25 -64290
rect 423 -64307 440 -64290
rect 672 -64307 689 -64290
rect 506 -64307 523 -64290
rect 257 -64307 274 -64290
rect 174 -64307 191 -64290
rect 755 -64307 772 -64290
rect 8 -64449 25 -64432
rect 423 -64449 440 -64432
rect 506 -64449 523 -64432
rect 257 -64449 274 -64432
rect 174 -64449 191 -64432
rect 755 -64449 772 -64432
rect 921 -64591 938 -64574
rect 8 -64591 25 -64574
rect 423 -64591 440 -64574
rect 506 -64591 523 -64574
rect 257 -64591 274 -64574
rect 174 -64591 191 -64574
rect 921 -64733 938 -64716
rect 8 -64733 25 -64716
rect 672 -64733 689 -64716
rect 423 -64733 440 -64716
rect 257 -64733 274 -64716
rect 174 -64733 191 -64716
rect 755 -64733 772 -64716
rect 921 -64875 938 -64858
rect 8 -64875 25 -64858
rect 423 -64875 440 -64858
rect 672 -64875 689 -64858
rect 257 -64875 274 -64858
rect 174 -64875 191 -64858
rect 755 -64875 772 -64858
rect 921 -65017 938 -65000
rect 8 -65017 25 -65000
rect 423 -65017 440 -65000
rect 257 -65017 274 -65000
rect 174 -65017 191 -65000
rect 921 -65159 938 -65142
rect 8 -65159 25 -65142
rect 672 -65159 689 -65142
rect 506 -65159 523 -65142
rect 257 -65159 274 -65142
rect 174 -65159 191 -65142
rect 755 -65159 772 -65142
rect 921 -65301 938 -65284
rect 8 -65301 25 -65284
rect 506 -65301 523 -65284
rect 257 -65301 274 -65284
rect 174 -65301 191 -65284
rect 755 -65301 772 -65284
rect 8 -65443 25 -65426
rect 506 -65443 523 -65426
rect 672 -65443 689 -65426
rect 257 -65443 274 -65426
rect 174 -65443 191 -65426
rect 755 -65443 772 -65426
rect 8 -65585 25 -65568
rect 672 -65585 689 -65568
rect 257 -65585 274 -65568
rect 174 -65585 191 -65568
rect 755 -65585 772 -65568
rect 8 -65727 25 -65710
rect 672 -65727 689 -65710
rect 506 -65727 523 -65710
rect 257 -65727 274 -65710
rect 174 -65727 191 -65710
rect 755 -65727 772 -65710
rect 423 -65727 440 -65710
rect 8 -65869 25 -65852
rect 423 -65869 440 -65852
rect 672 -65869 689 -65852
rect 506 -65869 523 -65852
rect 174 -65869 191 -65852
rect 755 -65869 772 -65852
rect 921 -66011 938 -65994
rect 8 -66011 25 -65994
rect 672 -66011 689 -65994
rect 423 -66011 440 -65994
rect 174 -66011 191 -65994
rect 755 -66011 772 -65994
rect 921 -66153 938 -66136
rect 8 -66153 25 -66136
rect 423 -66153 440 -66136
rect 174 -66153 191 -66136
rect 755 -66153 772 -66136
rect 921 -66295 938 -66278
rect 8 -66295 25 -66278
rect 672 -66295 689 -66278
rect 506 -66295 523 -66278
rect 174 -66295 191 -66278
rect 755 -66295 772 -66278
rect 921 -66437 938 -66420
rect 8 -66437 25 -66420
rect 506 -66437 523 -66420
rect 672 -66437 689 -66420
rect 174 -66437 191 -66420
rect 755 -66437 772 -66420
rect 921 -66579 938 -66562
rect 8 -66579 25 -66562
rect 672 -66579 689 -66562
rect 174 -66579 191 -66562
rect 8 -66721 25 -66704
rect 672 -66721 689 -66704
rect 506 -66721 523 -66704
rect 423 -66721 440 -66704
rect 257 -66721 274 -66704
rect 755 -66721 772 -66704
rect 921 -66863 938 -66846
rect 8 -66863 25 -66846
rect 423 -66863 440 -66846
rect 506 -66863 523 -66846
rect 672 -66863 689 -66846
rect 257 -66863 274 -66846
rect 755 -66863 772 -66846
rect 921 -67005 938 -66988
rect 8 -67005 25 -66988
rect 423 -67005 440 -66988
rect 257 -67005 274 -66988
rect 755 -67005 772 -66988
rect 921 -67147 938 -67130
rect 8 -67147 25 -67130
rect 672 -67147 689 -67130
rect 506 -67147 523 -67130
rect 257 -67147 274 -67130
rect 755 -67147 772 -67130
rect 921 -67289 938 -67272
rect 8 -67289 25 -67272
rect 672 -67289 689 -67272
rect 257 -67289 274 -67272
rect 755 -67289 772 -67272
rect 8 -67431 25 -67414
rect 672 -67431 689 -67414
rect 506 -67431 523 -67414
rect 423 -67431 440 -67414
rect 257 -67431 274 -67414
rect 755 -67431 772 -67414
rect 921 -67573 938 -67556
rect 8 -67573 25 -67556
rect 423 -67573 440 -67556
rect 506 -67573 523 -67556
rect 755 -67573 772 -67556
rect 921 -67715 938 -67698
rect 8 -67715 25 -67698
rect 423 -67715 440 -67698
rect 672 -67715 689 -67698
rect 755 -67715 772 -67698
rect 921 -67857 938 -67840
rect 8 -67857 25 -67840
rect 672 -67857 689 -67840
rect 506 -67857 523 -67840
rect 755 -67857 772 -67840
rect 921 -67999 938 -67982
rect 8 -67999 25 -67982
rect 672 -67999 689 -67982
rect 506 -67999 523 -67982
rect 755 -67999 772 -67982
rect 921 -68141 938 -68124
rect 8 -68141 25 -68124
rect 755 -68141 772 -68124
rect 921 -68283 938 -68266
rect 423 -68283 440 -68266
rect 672 -68283 689 -68266
rect 506 -68283 523 -68266
rect 257 -68283 274 -68266
rect 174 -68283 191 -68266
rect 921 -68425 938 -68408
rect 672 -68425 689 -68408
rect 423 -68425 440 -68408
rect 257 -68425 274 -68408
rect 174 -68425 191 -68408
rect 755 -68425 772 -68408
rect 921 -68567 938 -68550
rect 423 -68567 440 -68550
rect 672 -68567 689 -68550
rect 506 -68567 523 -68550
rect 257 -68567 274 -68550
rect 174 -68567 191 -68550
rect 921 -68709 938 -68692
rect 506 -68709 523 -68692
rect 672 -68709 689 -68692
rect 257 -68709 274 -68692
rect 174 -68709 191 -68692
rect 755 -68709 772 -68692
rect 921 -68851 938 -68834
rect 672 -68851 689 -68834
rect 257 -68851 274 -68834
rect 174 -68851 191 -68834
rect 921 -68993 938 -68976
rect 672 -68993 689 -68976
rect 506 -68993 523 -68976
rect 423 -68993 440 -68976
rect 174 -68993 191 -68976
rect 755 -68993 772 -68976
rect 921 -69135 938 -69118
rect 423 -69135 440 -69118
rect 506 -69135 523 -69118
rect 672 -69135 689 -69118
rect 174 -69135 191 -69118
rect 921 -69277 938 -69260
rect 423 -69277 440 -69260
rect 672 -69277 689 -69260
rect 506 -69277 523 -69260
rect 174 -69277 191 -69260
rect 755 -69277 772 -69260
rect 921 -69419 938 -69402
rect 672 -69419 689 -69402
rect 506 -69419 523 -69402
rect 174 -69419 191 -69402
rect 921 -69561 938 -69544
rect 672 -69561 689 -69544
rect 174 -69561 191 -69544
rect 755 -69561 772 -69544
rect 921 -69703 938 -69686
rect 257 -69703 274 -69686
rect 672 -69703 689 -69686
rect 506 -69703 523 -69686
rect 423 -69703 440 -69686
rect 174 -69703 191 -69686
rect 755 -69703 772 -69686
rect 921 -69845 938 -69828
rect 423 -69845 440 -69828
rect 506 -69845 523 -69828
rect 257 -69845 274 -69828
rect 755 -69845 772 -69828
rect 672 -69987 689 -69970
rect 423 -69987 440 -69970
rect 257 -69987 274 -69970
rect 755 -69987 772 -69970
rect 921 -70129 938 -70112
rect 423 -70129 440 -70112
rect 672 -70129 689 -70112
rect 257 -70129 274 -70112
rect 506 -70129 523 -70112
rect 755 -70129 772 -70112
rect 672 -70271 689 -70254
rect 506 -70271 523 -70254
rect 257 -70271 274 -70254
rect 755 -70271 772 -70254
rect 921 -70413 938 -70396
rect 672 -70413 689 -70396
rect 506 -70413 523 -70396
rect 257 -70413 274 -70396
rect 921 -70555 938 -70538
rect 257 -70555 274 -70538
rect 755 -70555 772 -70538
rect 921 -70697 938 -70680
rect 672 -70697 689 -70680
rect 506 -70697 523 -70680
rect 423 -70697 440 -70680
rect 755 -70697 772 -70680
rect 921 -70839 938 -70822
rect 423 -70839 440 -70822
rect 506 -70839 523 -70822
rect 755 -70839 772 -70822
rect 921 -70981 938 -70964
rect 672 -70981 689 -70964
rect 423 -70981 440 -70964
rect 755 -70981 772 -70964
rect 423 -71123 440 -71106
rect 672 -71123 689 -71106
rect 755 -71123 772 -71106
rect 921 -71265 938 -71248
rect 423 -71265 440 -71248
rect 672 -71265 689 -71248
rect 506 -71265 523 -71248
rect 755 -71265 772 -71248
rect 672 -71407 689 -71390
rect 506 -71407 523 -71390
rect 755 -71407 772 -71390
rect 921 -71549 938 -71532
rect 506 -71549 523 -71532
rect 755 -71549 772 -71532
rect 921 -71691 938 -71674
rect 672 -71691 689 -71674
rect 506 -71691 523 -71674
rect 755 -71691 772 -71674
rect 921 -71833 938 -71816
rect 672 -71833 689 -71816
rect 755 -71833 772 -71816
rect 921 -71975 938 -71958
rect 672 -71975 689 -71958
rect 755 -72117 772 -72100
rect 921 -72117 938 -72100
rect 921 -72259 938 -72242
rect 755 -72259 772 -72242
rect 921 -72401 938 -72384
<< poly >>
rect -51 -17 996 0
rect -67 -25 -34 8
rect -51 -88 996 -71
rect -67 -96 -34 -63
rect -51 -159 996 -142
rect -67 -167 -34 -134
rect -51 -230 996 -213
rect -67 -238 -34 -205
rect -51 -301 996 -284
rect -67 -309 -34 -276
rect -51 -372 996 -355
rect -67 -380 -34 -347
rect -51 -443 996 -426
rect -67 -451 -34 -418
rect -51 -514 996 -497
rect -67 -522 -34 -489
rect -51 -585 996 -568
rect -67 -593 -34 -560
rect -51 -656 996 -639
rect -67 -664 -34 -631
rect -51 -727 996 -710
rect -67 -735 -34 -702
rect -51 -798 996 -781
rect -67 -806 -34 -773
rect -51 -869 996 -852
rect -67 -877 -34 -844
rect -51 -940 996 -923
rect -67 -948 -34 -915
rect -51 -1011 996 -994
rect -67 -1019 -34 -986
rect -51 -1082 996 -1065
rect -67 -1090 -34 -1057
rect -51 -1153 996 -1136
rect -67 -1161 -34 -1128
rect -51 -1224 996 -1207
rect -67 -1232 -34 -1199
rect -51 -1295 996 -1278
rect -67 -1303 -34 -1270
rect -51 -1366 996 -1349
rect -67 -1374 -34 -1341
rect -51 -1437 996 -1420
rect -67 -1445 -34 -1412
rect -51 -1508 996 -1491
rect -67 -1516 -34 -1483
rect -51 -1579 996 -1562
rect -67 -1587 -34 -1554
rect -51 -1650 996 -1633
rect -67 -1658 -34 -1625
rect -51 -1721 996 -1704
rect -67 -1729 -34 -1696
rect -51 -1792 996 -1775
rect -67 -1800 -34 -1767
rect -51 -1863 996 -1846
rect -67 -1871 -34 -1838
rect -51 -1934 996 -1917
rect -67 -1942 -34 -1909
rect -51 -2005 996 -1988
rect -67 -2013 -34 -1980
rect -51 -2076 996 -2059
rect -67 -2084 -34 -2051
rect -51 -2147 996 -2130
rect -67 -2155 -34 -2122
rect -51 -2218 996 -2201
rect -67 -2226 -34 -2193
rect -51 -2289 996 -2272
rect -67 -2297 -34 -2264
rect -51 -2360 996 -2343
rect -67 -2368 -34 -2335
rect -51 -2431 996 -2414
rect -67 -2439 -34 -2406
rect -51 -2502 996 -2485
rect -67 -2510 -34 -2477
rect -51 -2573 996 -2556
rect -67 -2581 -34 -2548
rect -51 -2644 996 -2627
rect -67 -2652 -34 -2619
rect -51 -2715 996 -2698
rect -67 -2723 -34 -2690
rect -51 -2786 996 -2769
rect -67 -2794 -34 -2761
rect -51 -2857 996 -2840
rect -67 -2865 -34 -2832
rect -51 -2928 996 -2911
rect -67 -2936 -34 -2903
rect -51 -2999 996 -2982
rect -67 -3007 -34 -2974
rect -51 -3070 996 -3053
rect -67 -3078 -34 -3045
rect -51 -3141 996 -3124
rect -67 -3149 -34 -3116
rect -51 -3212 996 -3195
rect -67 -3220 -34 -3187
rect -51 -3283 996 -3266
rect -67 -3291 -34 -3258
rect -51 -3354 996 -3337
rect -67 -3362 -34 -3329
rect -51 -3425 996 -3408
rect -67 -3433 -34 -3400
rect -51 -3496 996 -3479
rect -67 -3504 -34 -3471
rect -51 -3567 996 -3550
rect -67 -3575 -34 -3542
rect -51 -3638 996 -3621
rect -67 -3646 -34 -3613
rect -51 -3709 996 -3692
rect -67 -3717 -34 -3684
rect -51 -3780 996 -3763
rect -67 -3788 -34 -3755
rect -51 -3851 996 -3834
rect -67 -3859 -34 -3826
rect -51 -3922 996 -3905
rect -67 -3930 -34 -3897
rect -51 -3993 996 -3976
rect -67 -4001 -34 -3968
rect -51 -4064 996 -4047
rect -67 -4072 -34 -4039
rect -51 -4135 996 -4118
rect -67 -4143 -34 -4110
rect -51 -4206 996 -4189
rect -67 -4214 -34 -4181
rect -51 -4277 996 -4260
rect -67 -4285 -34 -4252
rect -51 -4348 996 -4331
rect -67 -4356 -34 -4323
rect -51 -4419 996 -4402
rect -67 -4427 -34 -4394
rect -51 -4490 996 -4473
rect -67 -4498 -34 -4465
rect -51 -4561 996 -4544
rect -67 -4569 -34 -4536
rect -51 -4632 996 -4615
rect -67 -4640 -34 -4607
rect -51 -4703 996 -4686
rect -67 -4711 -34 -4678
rect -51 -4774 996 -4757
rect -67 -4782 -34 -4749
rect -51 -4845 996 -4828
rect -67 -4853 -34 -4820
rect -51 -4916 996 -4899
rect -67 -4924 -34 -4891
rect -51 -4987 996 -4970
rect -67 -4995 -34 -4962
rect -51 -5058 996 -5041
rect -67 -5066 -34 -5033
rect -51 -5129 996 -5112
rect -67 -5137 -34 -5104
rect -51 -5200 996 -5183
rect -67 -5208 -34 -5175
rect -51 -5271 996 -5254
rect -67 -5279 -34 -5246
rect -51 -5342 996 -5325
rect -67 -5350 -34 -5317
rect -51 -5413 996 -5396
rect -67 -5421 -34 -5388
rect -51 -5484 996 -5467
rect -67 -5492 -34 -5459
rect -51 -5555 996 -5538
rect -67 -5563 -34 -5530
rect -51 -5626 996 -5609
rect -67 -5634 -34 -5601
rect -51 -5697 996 -5680
rect -67 -5705 -34 -5672
rect -51 -5768 996 -5751
rect -67 -5776 -34 -5743
rect -51 -5839 996 -5822
rect -67 -5847 -34 -5814
rect -51 -5910 996 -5893
rect -67 -5918 -34 -5885
rect -51 -5981 996 -5964
rect -67 -5989 -34 -5956
rect -51 -6052 996 -6035
rect -67 -6060 -34 -6027
rect -51 -6123 996 -6106
rect -67 -6131 -34 -6098
rect -51 -6194 996 -6177
rect -67 -6202 -34 -6169
rect -51 -6265 996 -6248
rect -67 -6273 -34 -6240
rect -51 -6336 996 -6319
rect -67 -6344 -34 -6311
rect -51 -6407 996 -6390
rect -67 -6415 -34 -6382
rect -51 -6478 996 -6461
rect -67 -6486 -34 -6453
rect -51 -6549 996 -6532
rect -67 -6557 -34 -6524
rect -51 -6620 996 -6603
rect -67 -6628 -34 -6595
rect -51 -6691 996 -6674
rect -67 -6699 -34 -6666
rect -51 -6762 996 -6745
rect -67 -6770 -34 -6737
rect -51 -6833 996 -6816
rect -67 -6841 -34 -6808
rect -51 -6904 996 -6887
rect -67 -6912 -34 -6879
rect -51 -6975 996 -6958
rect -67 -6983 -34 -6950
rect -51 -7046 996 -7029
rect -67 -7054 -34 -7021
rect -51 -7117 996 -7100
rect -67 -7125 -34 -7092
rect -51 -7188 996 -7171
rect -67 -7196 -34 -7163
rect -51 -7259 996 -7242
rect -67 -7267 -34 -7234
rect -51 -7330 996 -7313
rect -67 -7338 -34 -7305
rect -51 -7401 996 -7384
rect -67 -7409 -34 -7376
rect -51 -7472 996 -7455
rect -67 -7480 -34 -7447
rect -51 -7543 996 -7526
rect -67 -7551 -34 -7518
rect -51 -7614 996 -7597
rect -67 -7622 -34 -7589
rect -51 -7685 996 -7668
rect -67 -7693 -34 -7660
rect -51 -7756 996 -7739
rect -67 -7764 -34 -7731
rect -51 -7827 996 -7810
rect -67 -7835 -34 -7802
rect -51 -7898 996 -7881
rect -67 -7906 -34 -7873
rect -51 -7969 996 -7952
rect -67 -7977 -34 -7944
rect -51 -8040 996 -8023
rect -67 -8048 -34 -8015
rect -51 -8111 996 -8094
rect -67 -8119 -34 -8086
rect -51 -8182 996 -8165
rect -67 -8190 -34 -8157
rect -51 -8253 996 -8236
rect -67 -8261 -34 -8228
rect -51 -8324 996 -8307
rect -67 -8332 -34 -8299
rect -51 -8395 996 -8378
rect -67 -8403 -34 -8370
rect -51 -8466 996 -8449
rect -67 -8474 -34 -8441
rect -51 -8537 996 -8520
rect -67 -8545 -34 -8512
rect -51 -8608 996 -8591
rect -67 -8616 -34 -8583
rect -51 -8679 996 -8662
rect -67 -8687 -34 -8654
rect -51 -8750 996 -8733
rect -67 -8758 -34 -8725
rect -51 -8821 996 -8804
rect -67 -8829 -34 -8796
rect -51 -8892 996 -8875
rect -67 -8900 -34 -8867
rect -51 -8963 996 -8946
rect -67 -8971 -34 -8938
rect -51 -9034 996 -9017
rect -67 -9042 -34 -9009
rect -51 -9105 996 -9088
rect -67 -9113 -34 -9080
rect -51 -9176 996 -9159
rect -67 -9184 -34 -9151
rect -51 -9247 996 -9230
rect -67 -9255 -34 -9222
rect -51 -9318 996 -9301
rect -67 -9326 -34 -9293
rect -51 -9389 996 -9372
rect -67 -9397 -34 -9364
rect -51 -9460 996 -9443
rect -67 -9468 -34 -9435
rect -51 -9531 996 -9514
rect -67 -9539 -34 -9506
rect -51 -9602 996 -9585
rect -67 -9610 -34 -9577
rect -51 -9673 996 -9656
rect -67 -9681 -34 -9648
rect -51 -9744 996 -9727
rect -67 -9752 -34 -9719
rect -51 -9815 996 -9798
rect -67 -9823 -34 -9790
rect -51 -9886 996 -9869
rect -67 -9894 -34 -9861
rect -51 -9957 996 -9940
rect -67 -9965 -34 -9932
rect -51 -10028 996 -10011
rect -67 -10036 -34 -10003
rect -51 -10099 996 -10082
rect -67 -10107 -34 -10074
rect -51 -10170 996 -10153
rect -67 -10178 -34 -10145
rect -51 -10241 996 -10224
rect -67 -10249 -34 -10216
rect -51 -10312 996 -10295
rect -67 -10320 -34 -10287
rect -51 -10383 996 -10366
rect -67 -10391 -34 -10358
rect -51 -10454 996 -10437
rect -67 -10462 -34 -10429
rect -51 -10525 996 -10508
rect -67 -10533 -34 -10500
rect -51 -10596 996 -10579
rect -67 -10604 -34 -10571
rect -51 -10667 996 -10650
rect -67 -10675 -34 -10642
rect -51 -10738 996 -10721
rect -67 -10746 -34 -10713
rect -51 -10809 996 -10792
rect -67 -10817 -34 -10784
rect -51 -10880 996 -10863
rect -67 -10888 -34 -10855
rect -51 -10951 996 -10934
rect -67 -10959 -34 -10926
rect -51 -11022 996 -11005
rect -67 -11030 -34 -10997
rect -51 -11093 996 -11076
rect -67 -11101 -34 -11068
rect -51 -11164 996 -11147
rect -67 -11172 -34 -11139
rect -51 -11235 996 -11218
rect -67 -11243 -34 -11210
rect -51 -11306 996 -11289
rect -67 -11314 -34 -11281
rect -51 -11377 996 -11360
rect -67 -11385 -34 -11352
rect -51 -11448 996 -11431
rect -67 -11456 -34 -11423
rect -51 -11519 996 -11502
rect -67 -11527 -34 -11494
rect -51 -11590 996 -11573
rect -67 -11598 -34 -11565
rect -51 -11661 996 -11644
rect -67 -11669 -34 -11636
rect -51 -11732 996 -11715
rect -67 -11740 -34 -11707
rect -51 -11803 996 -11786
rect -67 -11811 -34 -11778
rect -51 -11874 996 -11857
rect -67 -11882 -34 -11849
rect -51 -11945 996 -11928
rect -67 -11953 -34 -11920
rect -51 -12016 996 -11999
rect -67 -12024 -34 -11991
rect -51 -12087 996 -12070
rect -67 -12095 -34 -12062
rect -51 -12158 996 -12141
rect -67 -12166 -34 -12133
rect -51 -12229 996 -12212
rect -67 -12237 -34 -12204
rect -51 -12300 996 -12283
rect -67 -12308 -34 -12275
rect -51 -12371 996 -12354
rect -67 -12379 -34 -12346
rect -51 -12442 996 -12425
rect -67 -12450 -34 -12417
rect -51 -12513 996 -12496
rect -67 -12521 -34 -12488
rect -51 -12584 996 -12567
rect -67 -12592 -34 -12559
rect -51 -12655 996 -12638
rect -67 -12663 -34 -12630
rect -51 -12726 996 -12709
rect -67 -12734 -34 -12701
rect -51 -12797 996 -12780
rect -67 -12805 -34 -12772
rect -51 -12868 996 -12851
rect -67 -12876 -34 -12843
rect -51 -12939 996 -12922
rect -67 -12947 -34 -12914
rect -51 -13010 996 -12993
rect -67 -13018 -34 -12985
rect -51 -13081 996 -13064
rect -67 -13089 -34 -13056
rect -51 -13152 996 -13135
rect -67 -13160 -34 -13127
rect -51 -13223 996 -13206
rect -67 -13231 -34 -13198
rect -51 -13294 996 -13277
rect -67 -13302 -34 -13269
rect -51 -13365 996 -13348
rect -67 -13373 -34 -13340
rect -51 -13436 996 -13419
rect -67 -13444 -34 -13411
rect -51 -13507 996 -13490
rect -67 -13515 -34 -13482
rect -51 -13578 996 -13561
rect -67 -13586 -34 -13553
rect -51 -13649 996 -13632
rect -67 -13657 -34 -13624
rect -51 -13720 996 -13703
rect -67 -13728 -34 -13695
rect -51 -13791 996 -13774
rect -67 -13799 -34 -13766
rect -51 -13862 996 -13845
rect -67 -13870 -34 -13837
rect -51 -13933 996 -13916
rect -67 -13941 -34 -13908
rect -51 -14004 996 -13987
rect -67 -14012 -34 -13979
rect -51 -14075 996 -14058
rect -67 -14083 -34 -14050
rect -51 -14146 996 -14129
rect -67 -14154 -34 -14121
rect -51 -14217 996 -14200
rect -67 -14225 -34 -14192
rect -51 -14288 996 -14271
rect -67 -14296 -34 -14263
rect -51 -14359 996 -14342
rect -67 -14367 -34 -14334
rect -51 -14430 996 -14413
rect -67 -14438 -34 -14405
rect -51 -14501 996 -14484
rect -67 -14509 -34 -14476
rect -51 -14572 996 -14555
rect -67 -14580 -34 -14547
rect -51 -14643 996 -14626
rect -67 -14651 -34 -14618
rect -51 -14714 996 -14697
rect -67 -14722 -34 -14689
rect -51 -14785 996 -14768
rect -67 -14793 -34 -14760
rect -51 -14856 996 -14839
rect -67 -14864 -34 -14831
rect -51 -14927 996 -14910
rect -67 -14935 -34 -14902
rect -51 -14998 996 -14981
rect -67 -15006 -34 -14973
rect -51 -15069 996 -15052
rect -67 -15077 -34 -15044
rect -51 -15140 996 -15123
rect -67 -15148 -34 -15115
rect -51 -15211 996 -15194
rect -67 -15219 -34 -15186
rect -51 -15282 996 -15265
rect -67 -15290 -34 -15257
rect -51 -15353 996 -15336
rect -67 -15361 -34 -15328
rect -51 -15424 996 -15407
rect -67 -15432 -34 -15399
rect -51 -15495 996 -15478
rect -67 -15503 -34 -15470
rect -51 -15566 996 -15549
rect -67 -15574 -34 -15541
rect -51 -15637 996 -15620
rect -67 -15645 -34 -15612
rect -51 -15708 996 -15691
rect -67 -15716 -34 -15683
rect -51 -15779 996 -15762
rect -67 -15787 -34 -15754
rect -51 -15850 996 -15833
rect -67 -15858 -34 -15825
rect -51 -15921 996 -15904
rect -67 -15929 -34 -15896
rect -51 -15992 996 -15975
rect -67 -16000 -34 -15967
rect -51 -16063 996 -16046
rect -67 -16071 -34 -16038
rect -51 -16134 996 -16117
rect -67 -16142 -34 -16109
rect -51 -16205 996 -16188
rect -67 -16213 -34 -16180
rect -51 -16276 996 -16259
rect -67 -16284 -34 -16251
rect -51 -16347 996 -16330
rect -67 -16355 -34 -16322
rect -51 -16418 996 -16401
rect -67 -16426 -34 -16393
rect -51 -16489 996 -16472
rect -67 -16497 -34 -16464
rect -51 -16560 996 -16543
rect -67 -16568 -34 -16535
rect -51 -16631 996 -16614
rect -67 -16639 -34 -16606
rect -51 -16702 996 -16685
rect -67 -16710 -34 -16677
rect -51 -16773 996 -16756
rect -67 -16781 -34 -16748
rect -51 -16844 996 -16827
rect -67 -16852 -34 -16819
rect -51 -16915 996 -16898
rect -67 -16923 -34 -16890
rect -51 -16986 996 -16969
rect -67 -16994 -34 -16961
rect -51 -17057 996 -17040
rect -67 -17065 -34 -17032
rect -51 -17128 996 -17111
rect -67 -17136 -34 -17103
rect -51 -17199 996 -17182
rect -67 -17207 -34 -17174
rect -51 -17270 996 -17253
rect -67 -17278 -34 -17245
rect -51 -17341 996 -17324
rect -67 -17349 -34 -17316
rect -51 -17412 996 -17395
rect -67 -17420 -34 -17387
rect -51 -17483 996 -17466
rect -67 -17491 -34 -17458
rect -51 -17554 996 -17537
rect -67 -17562 -34 -17529
rect -51 -17625 996 -17608
rect -67 -17633 -34 -17600
rect -51 -17696 996 -17679
rect -67 -17704 -34 -17671
rect -51 -17767 996 -17750
rect -67 -17775 -34 -17742
rect -51 -17838 996 -17821
rect -67 -17846 -34 -17813
rect -51 -17909 996 -17892
rect -67 -17917 -34 -17884
rect -51 -17980 996 -17963
rect -67 -17988 -34 -17955
rect -51 -18051 996 -18034
rect -67 -18059 -34 -18026
rect -51 -18122 996 -18105
rect -67 -18130 -34 -18097
rect -51 -18193 996 -18176
rect -67 -18201 -34 -18168
rect -51 -18264 996 -18247
rect -67 -18272 -34 -18239
rect -51 -18335 996 -18318
rect -67 -18343 -34 -18310
rect -51 -18406 996 -18389
rect -67 -18414 -34 -18381
rect -51 -18477 996 -18460
rect -67 -18485 -34 -18452
rect -51 -18548 996 -18531
rect -67 -18556 -34 -18523
rect -51 -18619 996 -18602
rect -67 -18627 -34 -18594
rect -51 -18690 996 -18673
rect -67 -18698 -34 -18665
rect -51 -18761 996 -18744
rect -67 -18769 -34 -18736
rect -51 -18832 996 -18815
rect -67 -18840 -34 -18807
rect -51 -18903 996 -18886
rect -67 -18911 -34 -18878
rect -51 -18974 996 -18957
rect -67 -18982 -34 -18949
rect -51 -19045 996 -19028
rect -67 -19053 -34 -19020
rect -51 -19116 996 -19099
rect -67 -19124 -34 -19091
rect -51 -19187 996 -19170
rect -67 -19195 -34 -19162
rect -51 -19258 996 -19241
rect -67 -19266 -34 -19233
rect -51 -19329 996 -19312
rect -67 -19337 -34 -19304
rect -51 -19400 996 -19383
rect -67 -19408 -34 -19375
rect -51 -19471 996 -19454
rect -67 -19479 -34 -19446
rect -51 -19542 996 -19525
rect -67 -19550 -34 -19517
rect -51 -19613 996 -19596
rect -67 -19621 -34 -19588
rect -51 -19684 996 -19667
rect -67 -19692 -34 -19659
rect -51 -19755 996 -19738
rect -67 -19763 -34 -19730
rect -51 -19826 996 -19809
rect -67 -19834 -34 -19801
rect -51 -19897 996 -19880
rect -67 -19905 -34 -19872
rect -51 -19968 996 -19951
rect -67 -19976 -34 -19943
rect -51 -20039 996 -20022
rect -67 -20047 -34 -20014
rect -51 -20110 996 -20093
rect -67 -20118 -34 -20085
rect -51 -20181 996 -20164
rect -67 -20189 -34 -20156
rect -51 -20252 996 -20235
rect -67 -20260 -34 -20227
rect -51 -20323 996 -20306
rect -67 -20331 -34 -20298
rect -51 -20394 996 -20377
rect -67 -20402 -34 -20369
rect -51 -20465 996 -20448
rect -67 -20473 -34 -20440
rect -51 -20536 996 -20519
rect -67 -20544 -34 -20511
rect -51 -20607 996 -20590
rect -67 -20615 -34 -20582
rect -51 -20678 996 -20661
rect -67 -20686 -34 -20653
rect -51 -20749 996 -20732
rect -67 -20757 -34 -20724
rect -51 -20820 996 -20803
rect -67 -20828 -34 -20795
rect -51 -20891 996 -20874
rect -67 -20899 -34 -20866
rect -51 -20962 996 -20945
rect -67 -20970 -34 -20937
rect -51 -21033 996 -21016
rect -67 -21041 -34 -21008
rect -51 -21104 996 -21087
rect -67 -21112 -34 -21079
rect -51 -21175 996 -21158
rect -67 -21183 -34 -21150
rect -51 -21246 996 -21229
rect -67 -21254 -34 -21221
rect -51 -21317 996 -21300
rect -67 -21325 -34 -21292
rect -51 -21388 996 -21371
rect -67 -21396 -34 -21363
rect -51 -21459 996 -21442
rect -67 -21467 -34 -21434
rect -51 -21530 996 -21513
rect -67 -21538 -34 -21505
rect -51 -21601 996 -21584
rect -67 -21609 -34 -21576
rect -51 -21672 996 -21655
rect -67 -21680 -34 -21647
rect -51 -21743 996 -21726
rect -67 -21751 -34 -21718
rect -51 -21814 996 -21797
rect -67 -21822 -34 -21789
rect -51 -21885 996 -21868
rect -67 -21893 -34 -21860
rect -51 -21956 996 -21939
rect -67 -21964 -34 -21931
rect -51 -22027 996 -22010
rect -67 -22035 -34 -22002
rect -51 -22098 996 -22081
rect -67 -22106 -34 -22073
rect -51 -22169 996 -22152
rect -67 -22177 -34 -22144
rect -51 -22240 996 -22223
rect -67 -22248 -34 -22215
rect -51 -22311 996 -22294
rect -67 -22319 -34 -22286
rect -51 -22382 996 -22365
rect -67 -22390 -34 -22357
rect -51 -22453 996 -22436
rect -67 -22461 -34 -22428
rect -51 -22524 996 -22507
rect -67 -22532 -34 -22499
rect -51 -22595 996 -22578
rect -67 -22603 -34 -22570
rect -51 -22666 996 -22649
rect -67 -22674 -34 -22641
rect -51 -22737 996 -22720
rect -67 -22745 -34 -22712
rect -51 -22808 996 -22791
rect -67 -22816 -34 -22783
rect -51 -22879 996 -22862
rect -67 -22887 -34 -22854
rect -51 -22950 996 -22933
rect -67 -22958 -34 -22925
rect -51 -23021 996 -23004
rect -67 -23029 -34 -22996
rect -51 -23092 996 -23075
rect -67 -23100 -34 -23067
rect -51 -23163 996 -23146
rect -67 -23171 -34 -23138
rect -51 -23234 996 -23217
rect -67 -23242 -34 -23209
rect -51 -23305 996 -23288
rect -67 -23313 -34 -23280
rect -51 -23376 996 -23359
rect -67 -23384 -34 -23351
rect -51 -23447 996 -23430
rect -67 -23455 -34 -23422
rect -51 -23518 996 -23501
rect -67 -23526 -34 -23493
rect -51 -23589 996 -23572
rect -67 -23597 -34 -23564
rect -51 -23660 996 -23643
rect -67 -23668 -34 -23635
rect -51 -23731 996 -23714
rect -67 -23739 -34 -23706
rect -51 -23802 996 -23785
rect -67 -23810 -34 -23777
rect -51 -23873 996 -23856
rect -67 -23881 -34 -23848
rect -51 -23944 996 -23927
rect -67 -23952 -34 -23919
rect -51 -24015 996 -23998
rect -67 -24023 -34 -23990
rect -51 -24086 996 -24069
rect -67 -24094 -34 -24061
rect -51 -24157 996 -24140
rect -67 -24165 -34 -24132
rect -51 -24228 996 -24211
rect -67 -24236 -34 -24203
rect -51 -24299 996 -24282
rect -67 -24307 -34 -24274
rect -51 -24370 996 -24353
rect -67 -24378 -34 -24345
rect -51 -24441 996 -24424
rect -67 -24449 -34 -24416
rect -51 -24512 996 -24495
rect -67 -24520 -34 -24487
rect -51 -24583 996 -24566
rect -67 -24591 -34 -24558
rect -51 -24654 996 -24637
rect -67 -24662 -34 -24629
rect -51 -24725 996 -24708
rect -67 -24733 -34 -24700
rect -51 -24796 996 -24779
rect -67 -24804 -34 -24771
rect -51 -24867 996 -24850
rect -67 -24875 -34 -24842
rect -51 -24938 996 -24921
rect -67 -24946 -34 -24913
rect -51 -25009 996 -24992
rect -67 -25017 -34 -24984
rect -51 -25080 996 -25063
rect -67 -25088 -34 -25055
rect -51 -25151 996 -25134
rect -67 -25159 -34 -25126
rect -51 -25222 996 -25205
rect -67 -25230 -34 -25197
rect -51 -25293 996 -25276
rect -67 -25301 -34 -25268
rect -51 -25364 996 -25347
rect -67 -25372 -34 -25339
rect -51 -25435 996 -25418
rect -67 -25443 -34 -25410
rect -51 -25506 996 -25489
rect -67 -25514 -34 -25481
rect -51 -25577 996 -25560
rect -67 -25585 -34 -25552
rect -51 -25648 996 -25631
rect -67 -25656 -34 -25623
rect -51 -25719 996 -25702
rect -67 -25727 -34 -25694
rect -51 -25790 996 -25773
rect -67 -25798 -34 -25765
rect -51 -25861 996 -25844
rect -67 -25869 -34 -25836
rect -51 -25932 996 -25915
rect -67 -25940 -34 -25907
rect -51 -26003 996 -25986
rect -67 -26011 -34 -25978
rect -51 -26074 996 -26057
rect -67 -26082 -34 -26049
rect -51 -26145 996 -26128
rect -67 -26153 -34 -26120
rect -51 -26216 996 -26199
rect -67 -26224 -34 -26191
rect -51 -26287 996 -26270
rect -67 -26295 -34 -26262
rect -51 -26358 996 -26341
rect -67 -26366 -34 -26333
rect -51 -26429 996 -26412
rect -67 -26437 -34 -26404
rect -51 -26500 996 -26483
rect -67 -26508 -34 -26475
rect -51 -26571 996 -26554
rect -67 -26579 -34 -26546
rect -51 -26642 996 -26625
rect -67 -26650 -34 -26617
rect -51 -26713 996 -26696
rect -67 -26721 -34 -26688
rect -51 -26784 996 -26767
rect -67 -26792 -34 -26759
rect -51 -26855 996 -26838
rect -67 -26863 -34 -26830
rect -51 -26926 996 -26909
rect -67 -26934 -34 -26901
rect -51 -26997 996 -26980
rect -67 -27005 -34 -26972
rect -51 -27068 996 -27051
rect -67 -27076 -34 -27043
rect -51 -27139 996 -27122
rect -67 -27147 -34 -27114
rect -51 -27210 996 -27193
rect -67 -27218 -34 -27185
rect -51 -27281 996 -27264
rect -67 -27289 -34 -27256
rect -51 -27352 996 -27335
rect -67 -27360 -34 -27327
rect -51 -27423 996 -27406
rect -67 -27431 -34 -27398
rect -51 -27494 996 -27477
rect -67 -27502 -34 -27469
rect -51 -27565 996 -27548
rect -67 -27573 -34 -27540
rect -51 -27636 996 -27619
rect -67 -27644 -34 -27611
rect -51 -27707 996 -27690
rect -67 -27715 -34 -27682
rect -51 -27778 996 -27761
rect -67 -27786 -34 -27753
rect -51 -27849 996 -27832
rect -67 -27857 -34 -27824
rect -51 -27920 996 -27903
rect -67 -27928 -34 -27895
rect -51 -27991 996 -27974
rect -67 -27999 -34 -27966
rect -51 -28062 996 -28045
rect -67 -28070 -34 -28037
rect -51 -28133 996 -28116
rect -67 -28141 -34 -28108
rect -51 -28204 996 -28187
rect -67 -28212 -34 -28179
rect -51 -28275 996 -28258
rect -67 -28283 -34 -28250
rect -51 -28346 996 -28329
rect -67 -28354 -34 -28321
rect -51 -28417 996 -28400
rect -67 -28425 -34 -28392
rect -51 -28488 996 -28471
rect -67 -28496 -34 -28463
rect -51 -28559 996 -28542
rect -67 -28567 -34 -28534
rect -51 -28630 996 -28613
rect -67 -28638 -34 -28605
rect -51 -28701 996 -28684
rect -67 -28709 -34 -28676
rect -51 -28772 996 -28755
rect -67 -28780 -34 -28747
rect -51 -28843 996 -28826
rect -67 -28851 -34 -28818
rect -51 -28914 996 -28897
rect -67 -28922 -34 -28889
rect -51 -28985 996 -28968
rect -67 -28993 -34 -28960
rect -51 -29056 996 -29039
rect -67 -29064 -34 -29031
rect -51 -29127 996 -29110
rect -67 -29135 -34 -29102
rect -51 -29198 996 -29181
rect -67 -29206 -34 -29173
rect -51 -29269 996 -29252
rect -67 -29277 -34 -29244
rect -51 -29340 996 -29323
rect -67 -29348 -34 -29315
rect -51 -29411 996 -29394
rect -67 -29419 -34 -29386
rect -51 -29482 996 -29465
rect -67 -29490 -34 -29457
rect -51 -29553 996 -29536
rect -67 -29561 -34 -29528
rect -51 -29624 996 -29607
rect -67 -29632 -34 -29599
rect -51 -29695 996 -29678
rect -67 -29703 -34 -29670
rect -51 -29766 996 -29749
rect -67 -29774 -34 -29741
rect -51 -29837 996 -29820
rect -67 -29845 -34 -29812
rect -51 -29908 996 -29891
rect -67 -29916 -34 -29883
rect -51 -29979 996 -29962
rect -67 -29987 -34 -29954
rect -51 -30050 996 -30033
rect -67 -30058 -34 -30025
rect -51 -30121 996 -30104
rect -67 -30129 -34 -30096
rect -51 -30192 996 -30175
rect -67 -30200 -34 -30167
rect -51 -30263 996 -30246
rect -67 -30271 -34 -30238
rect -51 -30334 996 -30317
rect -67 -30342 -34 -30309
rect -51 -30405 996 -30388
rect -67 -30413 -34 -30380
rect -51 -30476 996 -30459
rect -67 -30484 -34 -30451
rect -51 -30547 996 -30530
rect -67 -30555 -34 -30522
rect -51 -30618 996 -30601
rect -67 -30626 -34 -30593
rect -51 -30689 996 -30672
rect -67 -30697 -34 -30664
rect -51 -30760 996 -30743
rect -67 -30768 -34 -30735
rect -51 -30831 996 -30814
rect -67 -30839 -34 -30806
rect -51 -30902 996 -30885
rect -67 -30910 -34 -30877
rect -51 -30973 996 -30956
rect -67 -30981 -34 -30948
rect -51 -31044 996 -31027
rect -67 -31052 -34 -31019
rect -51 -31115 996 -31098
rect -67 -31123 -34 -31090
rect -51 -31186 996 -31169
rect -67 -31194 -34 -31161
rect -51 -31257 996 -31240
rect -67 -31265 -34 -31232
rect -51 -31328 996 -31311
rect -67 -31336 -34 -31303
rect -51 -31399 996 -31382
rect -67 -31407 -34 -31374
rect -51 -31470 996 -31453
rect -67 -31478 -34 -31445
rect -51 -31541 996 -31524
rect -67 -31549 -34 -31516
rect -51 -31612 996 -31595
rect -67 -31620 -34 -31587
rect -51 -31683 996 -31666
rect -67 -31691 -34 -31658
rect -51 -31754 996 -31737
rect -67 -31762 -34 -31729
rect -51 -31825 996 -31808
rect -67 -31833 -34 -31800
rect -51 -31896 996 -31879
rect -67 -31904 -34 -31871
rect -51 -31967 996 -31950
rect -67 -31975 -34 -31942
rect -51 -32038 996 -32021
rect -67 -32046 -34 -32013
rect -51 -32109 996 -32092
rect -67 -32117 -34 -32084
rect -51 -32180 996 -32163
rect -67 -32188 -34 -32155
rect -51 -32251 996 -32234
rect -67 -32259 -34 -32226
rect -51 -32322 996 -32305
rect -67 -32330 -34 -32297
rect -51 -32393 996 -32376
rect -67 -32401 -34 -32368
rect -51 -32464 996 -32447
rect -67 -32472 -34 -32439
rect -51 -32535 996 -32518
rect -67 -32543 -34 -32510
rect -51 -32606 996 -32589
rect -67 -32614 -34 -32581
rect -51 -32677 996 -32660
rect -67 -32685 -34 -32652
rect -51 -32748 996 -32731
rect -67 -32756 -34 -32723
rect -51 -32819 996 -32802
rect -67 -32827 -34 -32794
rect -51 -32890 996 -32873
rect -67 -32898 -34 -32865
rect -51 -32961 996 -32944
rect -67 -32969 -34 -32936
rect -51 -33032 996 -33015
rect -67 -33040 -34 -33007
rect -51 -33103 996 -33086
rect -67 -33111 -34 -33078
rect -51 -33174 996 -33157
rect -67 -33182 -34 -33149
rect -51 -33245 996 -33228
rect -67 -33253 -34 -33220
rect -51 -33316 996 -33299
rect -67 -33324 -34 -33291
rect -51 -33387 996 -33370
rect -67 -33395 -34 -33362
rect -51 -33458 996 -33441
rect -67 -33466 -34 -33433
rect -51 -33529 996 -33512
rect -67 -33537 -34 -33504
rect -51 -33600 996 -33583
rect -67 -33608 -34 -33575
rect -51 -33671 996 -33654
rect -67 -33679 -34 -33646
rect -51 -33742 996 -33725
rect -67 -33750 -34 -33717
rect -51 -33813 996 -33796
rect -67 -33821 -34 -33788
rect -51 -33884 996 -33867
rect -67 -33892 -34 -33859
rect -51 -33955 996 -33938
rect -67 -33963 -34 -33930
rect -51 -34026 996 -34009
rect -67 -34034 -34 -34001
rect -51 -34097 996 -34080
rect -67 -34105 -34 -34072
rect -51 -34168 996 -34151
rect -67 -34176 -34 -34143
rect -51 -34239 996 -34222
rect -67 -34247 -34 -34214
rect -51 -34310 996 -34293
rect -67 -34318 -34 -34285
rect -51 -34381 996 -34364
rect -67 -34389 -34 -34356
rect -51 -34452 996 -34435
rect -67 -34460 -34 -34427
rect -51 -34523 996 -34506
rect -67 -34531 -34 -34498
rect -51 -34594 996 -34577
rect -67 -34602 -34 -34569
rect -51 -34665 996 -34648
rect -67 -34673 -34 -34640
rect -51 -34736 996 -34719
rect -67 -34744 -34 -34711
rect -51 -34807 996 -34790
rect -67 -34815 -34 -34782
rect -51 -34878 996 -34861
rect -67 -34886 -34 -34853
rect -51 -34949 996 -34932
rect -67 -34957 -34 -34924
rect -51 -35020 996 -35003
rect -67 -35028 -34 -34995
rect -51 -35091 996 -35074
rect -67 -35099 -34 -35066
rect -51 -35162 996 -35145
rect -67 -35170 -34 -35137
rect -51 -35233 996 -35216
rect -67 -35241 -34 -35208
rect -51 -35304 996 -35287
rect -67 -35312 -34 -35279
rect -51 -35375 996 -35358
rect -67 -35383 -34 -35350
rect -51 -35446 996 -35429
rect -67 -35454 -34 -35421
rect -51 -35517 996 -35500
rect -67 -35525 -34 -35492
rect -51 -35588 996 -35571
rect -67 -35596 -34 -35563
rect -51 -35659 996 -35642
rect -67 -35667 -34 -35634
rect -51 -35730 996 -35713
rect -67 -35738 -34 -35705
rect -51 -35801 996 -35784
rect -67 -35809 -34 -35776
rect -51 -35872 996 -35855
rect -67 -35880 -34 -35847
rect -51 -35943 996 -35926
rect -67 -35951 -34 -35918
rect -51 -36014 996 -35997
rect -67 -36022 -34 -35989
rect -51 -36085 996 -36068
rect -67 -36093 -34 -36060
rect -51 -36156 996 -36139
rect -67 -36164 -34 -36131
rect -51 -36227 996 -36210
rect -67 -36235 -34 -36202
rect -51 -36298 996 -36281
rect -67 -36306 -34 -36273
rect -51 -36369 996 -36352
rect -67 -36377 -34 -36344
rect -51 -36440 996 -36423
rect -67 -36448 -34 -36415
rect -51 -36511 996 -36494
rect -67 -36519 -34 -36486
rect -51 -36582 996 -36565
rect -67 -36590 -34 -36557
rect -51 -36653 996 -36636
rect -67 -36661 -34 -36628
rect -51 -36724 996 -36707
rect -67 -36732 -34 -36699
rect -51 -36795 996 -36778
rect -67 -36803 -34 -36770
rect -51 -36866 996 -36849
rect -67 -36874 -34 -36841
rect -51 -36937 996 -36920
rect -67 -36945 -34 -36912
rect -51 -37008 996 -36991
rect -67 -37016 -34 -36983
rect -51 -37079 996 -37062
rect -67 -37087 -34 -37054
rect -51 -37150 996 -37133
rect -67 -37158 -34 -37125
rect -51 -37221 996 -37204
rect -67 -37229 -34 -37196
rect -51 -37292 996 -37275
rect -67 -37300 -34 -37267
rect -51 -37363 996 -37346
rect -67 -37371 -34 -37338
rect -51 -37434 996 -37417
rect -67 -37442 -34 -37409
rect -51 -37505 996 -37488
rect -67 -37513 -34 -37480
rect -51 -37576 996 -37559
rect -67 -37584 -34 -37551
rect -51 -37647 996 -37630
rect -67 -37655 -34 -37622
rect -51 -37718 996 -37701
rect -67 -37726 -34 -37693
rect -51 -37789 996 -37772
rect -67 -37797 -34 -37764
rect -51 -37860 996 -37843
rect -67 -37868 -34 -37835
rect -51 -37931 996 -37914
rect -67 -37939 -34 -37906
rect -51 -38002 996 -37985
rect -67 -38010 -34 -37977
rect -51 -38073 996 -38056
rect -67 -38081 -34 -38048
rect -51 -38144 996 -38127
rect -67 -38152 -34 -38119
rect -51 -38215 996 -38198
rect -67 -38223 -34 -38190
rect -51 -38286 996 -38269
rect -67 -38294 -34 -38261
rect -51 -38357 996 -38340
rect -67 -38365 -34 -38332
rect -51 -38428 996 -38411
rect -67 -38436 -34 -38403
rect -51 -38499 996 -38482
rect -67 -38507 -34 -38474
rect -51 -38570 996 -38553
rect -67 -38578 -34 -38545
rect -51 -38641 996 -38624
rect -67 -38649 -34 -38616
rect -51 -38712 996 -38695
rect -67 -38720 -34 -38687
rect -51 -38783 996 -38766
rect -67 -38791 -34 -38758
rect -51 -38854 996 -38837
rect -67 -38862 -34 -38829
rect -51 -38925 996 -38908
rect -67 -38933 -34 -38900
rect -51 -38996 996 -38979
rect -67 -39004 -34 -38971
rect -51 -39067 996 -39050
rect -67 -39075 -34 -39042
rect -51 -39138 996 -39121
rect -67 -39146 -34 -39113
rect -51 -39209 996 -39192
rect -67 -39217 -34 -39184
rect -51 -39280 996 -39263
rect -67 -39288 -34 -39255
rect -51 -39351 996 -39334
rect -67 -39359 -34 -39326
rect -51 -39422 996 -39405
rect -67 -39430 -34 -39397
rect -51 -39493 996 -39476
rect -67 -39501 -34 -39468
rect -51 -39564 996 -39547
rect -67 -39572 -34 -39539
rect -51 -39635 996 -39618
rect -67 -39643 -34 -39610
rect -51 -39706 996 -39689
rect -67 -39714 -34 -39681
rect -51 -39777 996 -39760
rect -67 -39785 -34 -39752
rect -51 -39848 996 -39831
rect -67 -39856 -34 -39823
rect -51 -39919 996 -39902
rect -67 -39927 -34 -39894
rect -51 -39990 996 -39973
rect -67 -39998 -34 -39965
rect -51 -40061 996 -40044
rect -67 -40069 -34 -40036
rect -51 -40132 996 -40115
rect -67 -40140 -34 -40107
rect -51 -40203 996 -40186
rect -67 -40211 -34 -40178
rect -51 -40274 996 -40257
rect -67 -40282 -34 -40249
rect -51 -40345 996 -40328
rect -67 -40353 -34 -40320
rect -51 -40416 996 -40399
rect -67 -40424 -34 -40391
rect -51 -40487 996 -40470
rect -67 -40495 -34 -40462
rect -51 -40558 996 -40541
rect -67 -40566 -34 -40533
rect -51 -40629 996 -40612
rect -67 -40637 -34 -40604
rect -51 -40700 996 -40683
rect -67 -40708 -34 -40675
rect -51 -40771 996 -40754
rect -67 -40779 -34 -40746
rect -51 -40842 996 -40825
rect -67 -40850 -34 -40817
rect -51 -40913 996 -40896
rect -67 -40921 -34 -40888
rect -51 -40984 996 -40967
rect -67 -40992 -34 -40959
rect -51 -41055 996 -41038
rect -67 -41063 -34 -41030
rect -51 -41126 996 -41109
rect -67 -41134 -34 -41101
rect -51 -41197 996 -41180
rect -67 -41205 -34 -41172
rect -51 -41268 996 -41251
rect -67 -41276 -34 -41243
rect -51 -41339 996 -41322
rect -67 -41347 -34 -41314
rect -51 -41410 996 -41393
rect -67 -41418 -34 -41385
rect -51 -41481 996 -41464
rect -67 -41489 -34 -41456
rect -51 -41552 996 -41535
rect -67 -41560 -34 -41527
rect -51 -41623 996 -41606
rect -67 -41631 -34 -41598
rect -51 -41694 996 -41677
rect -67 -41702 -34 -41669
rect -51 -41765 996 -41748
rect -67 -41773 -34 -41740
rect -51 -41836 996 -41819
rect -67 -41844 -34 -41811
rect -51 -41907 996 -41890
rect -67 -41915 -34 -41882
rect -51 -41978 996 -41961
rect -67 -41986 -34 -41953
rect -51 -42049 996 -42032
rect -67 -42057 -34 -42024
rect -51 -42120 996 -42103
rect -67 -42128 -34 -42095
rect -51 -42191 996 -42174
rect -67 -42199 -34 -42166
rect -51 -42262 996 -42245
rect -67 -42270 -34 -42237
rect -51 -42333 996 -42316
rect -67 -42341 -34 -42308
rect -51 -42404 996 -42387
rect -67 -42412 -34 -42379
rect -51 -42475 996 -42458
rect -67 -42483 -34 -42450
rect -51 -42546 996 -42529
rect -67 -42554 -34 -42521
rect -51 -42617 996 -42600
rect -67 -42625 -34 -42592
rect -51 -42688 996 -42671
rect -67 -42696 -34 -42663
rect -51 -42759 996 -42742
rect -67 -42767 -34 -42734
rect -51 -42830 996 -42813
rect -67 -42838 -34 -42805
rect -51 -42901 996 -42884
rect -67 -42909 -34 -42876
rect -51 -42972 996 -42955
rect -67 -42980 -34 -42947
rect -51 -43043 996 -43026
rect -67 -43051 -34 -43018
rect -51 -43114 996 -43097
rect -67 -43122 -34 -43089
rect -51 -43185 996 -43168
rect -67 -43193 -34 -43160
rect -51 -43256 996 -43239
rect -67 -43264 -34 -43231
rect -51 -43327 996 -43310
rect -67 -43335 -34 -43302
rect -51 -43398 996 -43381
rect -67 -43406 -34 -43373
rect -51 -43469 996 -43452
rect -67 -43477 -34 -43444
rect -51 -43540 996 -43523
rect -67 -43548 -34 -43515
rect -51 -43611 996 -43594
rect -67 -43619 -34 -43586
rect -51 -43682 996 -43665
rect -67 -43690 -34 -43657
rect -51 -43753 996 -43736
rect -67 -43761 -34 -43728
rect -51 -43824 996 -43807
rect -67 -43832 -34 -43799
rect -51 -43895 996 -43878
rect -67 -43903 -34 -43870
rect -51 -43966 996 -43949
rect -67 -43974 -34 -43941
rect -51 -44037 996 -44020
rect -67 -44045 -34 -44012
rect -51 -44108 996 -44091
rect -67 -44116 -34 -44083
rect -51 -44179 996 -44162
rect -67 -44187 -34 -44154
rect -51 -44250 996 -44233
rect -67 -44258 -34 -44225
rect -51 -44321 996 -44304
rect -67 -44329 -34 -44296
rect -51 -44392 996 -44375
rect -67 -44400 -34 -44367
rect -51 -44463 996 -44446
rect -67 -44471 -34 -44438
rect -51 -44534 996 -44517
rect -67 -44542 -34 -44509
rect -51 -44605 996 -44588
rect -67 -44613 -34 -44580
rect -51 -44676 996 -44659
rect -67 -44684 -34 -44651
rect -51 -44747 996 -44730
rect -67 -44755 -34 -44722
rect -51 -44818 996 -44801
rect -67 -44826 -34 -44793
rect -51 -44889 996 -44872
rect -67 -44897 -34 -44864
rect -51 -44960 996 -44943
rect -67 -44968 -34 -44935
rect -51 -45031 996 -45014
rect -67 -45039 -34 -45006
rect -51 -45102 996 -45085
rect -67 -45110 -34 -45077
rect -51 -45173 996 -45156
rect -67 -45181 -34 -45148
rect -51 -45244 996 -45227
rect -67 -45252 -34 -45219
rect -51 -45315 996 -45298
rect -67 -45323 -34 -45290
rect -51 -45386 996 -45369
rect -67 -45394 -34 -45361
rect -51 -45457 996 -45440
rect -67 -45465 -34 -45432
rect -51 -45528 996 -45511
rect -67 -45536 -34 -45503
rect -51 -45599 996 -45582
rect -67 -45607 -34 -45574
rect -51 -45670 996 -45653
rect -67 -45678 -34 -45645
rect -51 -45741 996 -45724
rect -67 -45749 -34 -45716
rect -51 -45812 996 -45795
rect -67 -45820 -34 -45787
rect -51 -45883 996 -45866
rect -67 -45891 -34 -45858
rect -51 -45954 996 -45937
rect -67 -45962 -34 -45929
rect -51 -46025 996 -46008
rect -67 -46033 -34 -46000
rect -51 -46096 996 -46079
rect -67 -46104 -34 -46071
rect -51 -46167 996 -46150
rect -67 -46175 -34 -46142
rect -51 -46238 996 -46221
rect -67 -46246 -34 -46213
rect -51 -46309 996 -46292
rect -67 -46317 -34 -46284
rect -51 -46380 996 -46363
rect -67 -46388 -34 -46355
rect -51 -46451 996 -46434
rect -67 -46459 -34 -46426
rect -51 -46522 996 -46505
rect -67 -46530 -34 -46497
rect -51 -46593 996 -46576
rect -67 -46601 -34 -46568
rect -51 -46664 996 -46647
rect -67 -46672 -34 -46639
rect -51 -46735 996 -46718
rect -67 -46743 -34 -46710
rect -51 -46806 996 -46789
rect -67 -46814 -34 -46781
rect -51 -46877 996 -46860
rect -67 -46885 -34 -46852
rect -51 -46948 996 -46931
rect -67 -46956 -34 -46923
rect -51 -47019 996 -47002
rect -67 -47027 -34 -46994
rect -51 -47090 996 -47073
rect -67 -47098 -34 -47065
rect -51 -47161 996 -47144
rect -67 -47169 -34 -47136
rect -51 -47232 996 -47215
rect -67 -47240 -34 -47207
rect -51 -47303 996 -47286
rect -67 -47311 -34 -47278
rect -51 -47374 996 -47357
rect -67 -47382 -34 -47349
rect -51 -47445 996 -47428
rect -67 -47453 -34 -47420
rect -51 -47516 996 -47499
rect -67 -47524 -34 -47491
rect -51 -47587 996 -47570
rect -67 -47595 -34 -47562
rect -51 -47658 996 -47641
rect -67 -47666 -34 -47633
rect -51 -47729 996 -47712
rect -67 -47737 -34 -47704
rect -51 -47800 996 -47783
rect -67 -47808 -34 -47775
rect -51 -47871 996 -47854
rect -67 -47879 -34 -47846
rect -51 -47942 996 -47925
rect -67 -47950 -34 -47917
rect -51 -48013 996 -47996
rect -67 -48021 -34 -47988
rect -51 -48084 996 -48067
rect -67 -48092 -34 -48059
rect -51 -48155 996 -48138
rect -67 -48163 -34 -48130
rect -51 -48226 996 -48209
rect -67 -48234 -34 -48201
rect -51 -48297 996 -48280
rect -67 -48305 -34 -48272
rect -51 -48368 996 -48351
rect -67 -48376 -34 -48343
rect -51 -48439 996 -48422
rect -67 -48447 -34 -48414
rect -51 -48510 996 -48493
rect -67 -48518 -34 -48485
rect -51 -48581 996 -48564
rect -67 -48589 -34 -48556
rect -51 -48652 996 -48635
rect -67 -48660 -34 -48627
rect -51 -48723 996 -48706
rect -67 -48731 -34 -48698
rect -51 -48794 996 -48777
rect -67 -48802 -34 -48769
rect -51 -48865 996 -48848
rect -67 -48873 -34 -48840
rect -51 -48936 996 -48919
rect -67 -48944 -34 -48911
rect -51 -49007 996 -48990
rect -67 -49015 -34 -48982
rect -51 -49078 996 -49061
rect -67 -49086 -34 -49053
rect -51 -49149 996 -49132
rect -67 -49157 -34 -49124
rect -51 -49220 996 -49203
rect -67 -49228 -34 -49195
rect -51 -49291 996 -49274
rect -67 -49299 -34 -49266
rect -51 -49362 996 -49345
rect -67 -49370 -34 -49337
rect -51 -49433 996 -49416
rect -67 -49441 -34 -49408
rect -51 -49504 996 -49487
rect -67 -49512 -34 -49479
rect -51 -49575 996 -49558
rect -67 -49583 -34 -49550
rect -51 -49646 996 -49629
rect -67 -49654 -34 -49621
rect -51 -49717 996 -49700
rect -67 -49725 -34 -49692
rect -51 -49788 996 -49771
rect -67 -49796 -34 -49763
rect -51 -49859 996 -49842
rect -67 -49867 -34 -49834
rect -51 -49930 996 -49913
rect -67 -49938 -34 -49905
rect -51 -50001 996 -49984
rect -67 -50009 -34 -49976
rect -51 -50072 996 -50055
rect -67 -50080 -34 -50047
rect -51 -50143 996 -50126
rect -67 -50151 -34 -50118
rect -51 -50214 996 -50197
rect -67 -50222 -34 -50189
rect -51 -50285 996 -50268
rect -67 -50293 -34 -50260
rect -51 -50356 996 -50339
rect -67 -50364 -34 -50331
rect -51 -50427 996 -50410
rect -67 -50435 -34 -50402
rect -51 -50498 996 -50481
rect -67 -50506 -34 -50473
rect -51 -50569 996 -50552
rect -67 -50577 -34 -50544
rect -51 -50640 996 -50623
rect -67 -50648 -34 -50615
rect -51 -50711 996 -50694
rect -67 -50719 -34 -50686
rect -51 -50782 996 -50765
rect -67 -50790 -34 -50757
rect -51 -50853 996 -50836
rect -67 -50861 -34 -50828
rect -51 -50924 996 -50907
rect -67 -50932 -34 -50899
rect -51 -50995 996 -50978
rect -67 -51003 -34 -50970
rect -51 -51066 996 -51049
rect -67 -51074 -34 -51041
rect -51 -51137 996 -51120
rect -67 -51145 -34 -51112
rect -51 -51208 996 -51191
rect -67 -51216 -34 -51183
rect -51 -51279 996 -51262
rect -67 -51287 -34 -51254
rect -51 -51350 996 -51333
rect -67 -51358 -34 -51325
rect -51 -51421 996 -51404
rect -67 -51429 -34 -51396
rect -51 -51492 996 -51475
rect -67 -51500 -34 -51467
rect -51 -51563 996 -51546
rect -67 -51571 -34 -51538
rect -51 -51634 996 -51617
rect -67 -51642 -34 -51609
rect -51 -51705 996 -51688
rect -67 -51713 -34 -51680
rect -51 -51776 996 -51759
rect -67 -51784 -34 -51751
rect -51 -51847 996 -51830
rect -67 -51855 -34 -51822
rect -51 -51918 996 -51901
rect -67 -51926 -34 -51893
rect -51 -51989 996 -51972
rect -67 -51997 -34 -51964
rect -51 -52060 996 -52043
rect -67 -52068 -34 -52035
rect -51 -52131 996 -52114
rect -67 -52139 -34 -52106
rect -51 -52202 996 -52185
rect -67 -52210 -34 -52177
rect -51 -52273 996 -52256
rect -67 -52281 -34 -52248
rect -51 -52344 996 -52327
rect -67 -52352 -34 -52319
rect -51 -52415 996 -52398
rect -67 -52423 -34 -52390
rect -51 -52486 996 -52469
rect -67 -52494 -34 -52461
rect -51 -52557 996 -52540
rect -67 -52565 -34 -52532
rect -51 -52628 996 -52611
rect -67 -52636 -34 -52603
rect -51 -52699 996 -52682
rect -67 -52707 -34 -52674
rect -51 -52770 996 -52753
rect -67 -52778 -34 -52745
rect -51 -52841 996 -52824
rect -67 -52849 -34 -52816
rect -51 -52912 996 -52895
rect -67 -52920 -34 -52887
rect -51 -52983 996 -52966
rect -67 -52991 -34 -52958
rect -51 -53054 996 -53037
rect -67 -53062 -34 -53029
rect -51 -53125 996 -53108
rect -67 -53133 -34 -53100
rect -51 -53196 996 -53179
rect -67 -53204 -34 -53171
rect -51 -53267 996 -53250
rect -67 -53275 -34 -53242
rect -51 -53338 996 -53321
rect -67 -53346 -34 -53313
rect -51 -53409 996 -53392
rect -67 -53417 -34 -53384
rect -51 -53480 996 -53463
rect -67 -53488 -34 -53455
rect -51 -53551 996 -53534
rect -67 -53559 -34 -53526
rect -51 -53622 996 -53605
rect -67 -53630 -34 -53597
rect -51 -53693 996 -53676
rect -67 -53701 -34 -53668
rect -51 -53764 996 -53747
rect -67 -53772 -34 -53739
rect -51 -53835 996 -53818
rect -67 -53843 -34 -53810
rect -51 -53906 996 -53889
rect -67 -53914 -34 -53881
rect -51 -53977 996 -53960
rect -67 -53985 -34 -53952
rect -51 -54048 996 -54031
rect -67 -54056 -34 -54023
rect -51 -54119 996 -54102
rect -67 -54127 -34 -54094
rect -51 -54190 996 -54173
rect -67 -54198 -34 -54165
rect -51 -54261 996 -54244
rect -67 -54269 -34 -54236
rect -51 -54332 996 -54315
rect -67 -54340 -34 -54307
rect -51 -54403 996 -54386
rect -67 -54411 -34 -54378
rect -51 -54474 996 -54457
rect -67 -54482 -34 -54449
rect -51 -54545 996 -54528
rect -67 -54553 -34 -54520
rect -51 -54616 996 -54599
rect -67 -54624 -34 -54591
rect -51 -54687 996 -54670
rect -67 -54695 -34 -54662
rect -51 -54758 996 -54741
rect -67 -54766 -34 -54733
rect -51 -54829 996 -54812
rect -67 -54837 -34 -54804
rect -51 -54900 996 -54883
rect -67 -54908 -34 -54875
rect -51 -54971 996 -54954
rect -67 -54979 -34 -54946
rect -51 -55042 996 -55025
rect -67 -55050 -34 -55017
rect -51 -55113 996 -55096
rect -67 -55121 -34 -55088
rect -51 -55184 996 -55167
rect -67 -55192 -34 -55159
rect -51 -55255 996 -55238
rect -67 -55263 -34 -55230
rect -51 -55326 996 -55309
rect -67 -55334 -34 -55301
rect -51 -55397 996 -55380
rect -67 -55405 -34 -55372
rect -51 -55468 996 -55451
rect -67 -55476 -34 -55443
rect -51 -55539 996 -55522
rect -67 -55547 -34 -55514
rect -51 -55610 996 -55593
rect -67 -55618 -34 -55585
rect -51 -55681 996 -55664
rect -67 -55689 -34 -55656
rect -51 -55752 996 -55735
rect -67 -55760 -34 -55727
rect -51 -55823 996 -55806
rect -67 -55831 -34 -55798
rect -51 -55894 996 -55877
rect -67 -55902 -34 -55869
rect -51 -55965 996 -55948
rect -67 -55973 -34 -55940
rect -51 -56036 996 -56019
rect -67 -56044 -34 -56011
rect -51 -56107 996 -56090
rect -67 -56115 -34 -56082
rect -51 -56178 996 -56161
rect -67 -56186 -34 -56153
rect -51 -56249 996 -56232
rect -67 -56257 -34 -56224
rect -51 -56320 996 -56303
rect -67 -56328 -34 -56295
rect -51 -56391 996 -56374
rect -67 -56399 -34 -56366
rect -51 -56462 996 -56445
rect -67 -56470 -34 -56437
rect -51 -56533 996 -56516
rect -67 -56541 -34 -56508
rect -51 -56604 996 -56587
rect -67 -56612 -34 -56579
rect -51 -56675 996 -56658
rect -67 -56683 -34 -56650
rect -51 -56746 996 -56729
rect -67 -56754 -34 -56721
rect -51 -56817 996 -56800
rect -67 -56825 -34 -56792
rect -51 -56888 996 -56871
rect -67 -56896 -34 -56863
rect -51 -56959 996 -56942
rect -67 -56967 -34 -56934
rect -51 -57030 996 -57013
rect -67 -57038 -34 -57005
rect -51 -57101 996 -57084
rect -67 -57109 -34 -57076
rect -51 -57172 996 -57155
rect -67 -57180 -34 -57147
rect -51 -57243 996 -57226
rect -67 -57251 -34 -57218
rect -51 -57314 996 -57297
rect -67 -57322 -34 -57289
rect -51 -57385 996 -57368
rect -67 -57393 -34 -57360
rect -51 -57456 996 -57439
rect -67 -57464 -34 -57431
rect -51 -57527 996 -57510
rect -67 -57535 -34 -57502
rect -51 -57598 996 -57581
rect -67 -57606 -34 -57573
rect -51 -57669 996 -57652
rect -67 -57677 -34 -57644
rect -51 -57740 996 -57723
rect -67 -57748 -34 -57715
rect -51 -57811 996 -57794
rect -67 -57819 -34 -57786
rect -51 -57882 996 -57865
rect -67 -57890 -34 -57857
rect -51 -57953 996 -57936
rect -67 -57961 -34 -57928
rect -51 -58024 996 -58007
rect -67 -58032 -34 -57999
rect -51 -58095 996 -58078
rect -67 -58103 -34 -58070
rect -51 -58166 996 -58149
rect -67 -58174 -34 -58141
rect -51 -58237 996 -58220
rect -67 -58245 -34 -58212
rect -51 -58308 996 -58291
rect -67 -58316 -34 -58283
rect -51 -58379 996 -58362
rect -67 -58387 -34 -58354
rect -51 -58450 996 -58433
rect -67 -58458 -34 -58425
rect -51 -58521 996 -58504
rect -67 -58529 -34 -58496
rect -51 -58592 996 -58575
rect -67 -58600 -34 -58567
rect -51 -58663 996 -58646
rect -67 -58671 -34 -58638
rect -51 -58734 996 -58717
rect -67 -58742 -34 -58709
rect -51 -58805 996 -58788
rect -67 -58813 -34 -58780
rect -51 -58876 996 -58859
rect -67 -58884 -34 -58851
rect -51 -58947 996 -58930
rect -67 -58955 -34 -58922
rect -51 -59018 996 -59001
rect -67 -59026 -34 -58993
rect -51 -59089 996 -59072
rect -67 -59097 -34 -59064
rect -51 -59160 996 -59143
rect -67 -59168 -34 -59135
rect -51 -59231 996 -59214
rect -67 -59239 -34 -59206
rect -51 -59302 996 -59285
rect -67 -59310 -34 -59277
rect -51 -59373 996 -59356
rect -67 -59381 -34 -59348
rect -51 -59444 996 -59427
rect -67 -59452 -34 -59419
rect -51 -59515 996 -59498
rect -67 -59523 -34 -59490
rect -51 -59586 996 -59569
rect -67 -59594 -34 -59561
rect -51 -59657 996 -59640
rect -67 -59665 -34 -59632
rect -51 -59728 996 -59711
rect -67 -59736 -34 -59703
rect -51 -59799 996 -59782
rect -67 -59807 -34 -59774
rect -51 -59870 996 -59853
rect -67 -59878 -34 -59845
rect -51 -59941 996 -59924
rect -67 -59949 -34 -59916
rect -51 -60012 996 -59995
rect -67 -60020 -34 -59987
rect -51 -60083 996 -60066
rect -67 -60091 -34 -60058
rect -51 -60154 996 -60137
rect -67 -60162 -34 -60129
rect -51 -60225 996 -60208
rect -67 -60233 -34 -60200
rect -51 -60296 996 -60279
rect -67 -60304 -34 -60271
rect -51 -60367 996 -60350
rect -67 -60375 -34 -60342
rect -51 -60438 996 -60421
rect -67 -60446 -34 -60413
rect -51 -60509 996 -60492
rect -67 -60517 -34 -60484
rect -51 -60580 996 -60563
rect -67 -60588 -34 -60555
rect -51 -60651 996 -60634
rect -67 -60659 -34 -60626
rect -51 -60722 996 -60705
rect -67 -60730 -34 -60697
rect -51 -60793 996 -60776
rect -67 -60801 -34 -60768
rect -51 -60864 996 -60847
rect -67 -60872 -34 -60839
rect -51 -60935 996 -60918
rect -67 -60943 -34 -60910
rect -51 -61006 996 -60989
rect -67 -61014 -34 -60981
rect -51 -61077 996 -61060
rect -67 -61085 -34 -61052
rect -51 -61148 996 -61131
rect -67 -61156 -34 -61123
rect -51 -61219 996 -61202
rect -67 -61227 -34 -61194
rect -51 -61290 996 -61273
rect -67 -61298 -34 -61265
rect -51 -61361 996 -61344
rect -67 -61369 -34 -61336
rect -51 -61432 996 -61415
rect -67 -61440 -34 -61407
rect -51 -61503 996 -61486
rect -67 -61511 -34 -61478
rect -51 -61574 996 -61557
rect -67 -61582 -34 -61549
rect -51 -61645 996 -61628
rect -67 -61653 -34 -61620
rect -51 -61716 996 -61699
rect -67 -61724 -34 -61691
rect -51 -61787 996 -61770
rect -67 -61795 -34 -61762
rect -51 -61858 996 -61841
rect -67 -61866 -34 -61833
rect -51 -61929 996 -61912
rect -67 -61937 -34 -61904
rect -51 -62000 996 -61983
rect -67 -62008 -34 -61975
rect -51 -62071 996 -62054
rect -67 -62079 -34 -62046
rect -51 -62142 996 -62125
rect -67 -62150 -34 -62117
rect -51 -62213 996 -62196
rect -67 -62221 -34 -62188
rect -51 -62284 996 -62267
rect -67 -62292 -34 -62259
rect -51 -62355 996 -62338
rect -67 -62363 -34 -62330
rect -51 -62426 996 -62409
rect -67 -62434 -34 -62401
rect -51 -62497 996 -62480
rect -67 -62505 -34 -62472
rect -51 -62568 996 -62551
rect -67 -62576 -34 -62543
rect -51 -62639 996 -62622
rect -67 -62647 -34 -62614
rect -51 -62710 996 -62693
rect -67 -62718 -34 -62685
rect -51 -62781 996 -62764
rect -67 -62789 -34 -62756
rect -51 -62852 996 -62835
rect -67 -62860 -34 -62827
rect -51 -62923 996 -62906
rect -67 -62931 -34 -62898
rect -51 -62994 996 -62977
rect -67 -63002 -34 -62969
rect -51 -63065 996 -63048
rect -67 -63073 -34 -63040
rect -51 -63136 996 -63119
rect -67 -63144 -34 -63111
rect -51 -63207 996 -63190
rect -67 -63215 -34 -63182
rect -51 -63278 996 -63261
rect -67 -63286 -34 -63253
rect -51 -63349 996 -63332
rect -67 -63357 -34 -63324
rect -51 -63420 996 -63403
rect -67 -63428 -34 -63395
rect -51 -63491 996 -63474
rect -67 -63499 -34 -63466
rect -51 -63562 996 -63545
rect -67 -63570 -34 -63537
rect -51 -63633 996 -63616
rect -67 -63641 -34 -63608
rect -51 -63704 996 -63687
rect -67 -63712 -34 -63679
rect -51 -63775 996 -63758
rect -67 -63783 -34 -63750
rect -51 -63846 996 -63829
rect -67 -63854 -34 -63821
rect -51 -63917 996 -63900
rect -67 -63925 -34 -63892
rect -51 -63988 996 -63971
rect -67 -63996 -34 -63963
rect -51 -64059 996 -64042
rect -67 -64067 -34 -64034
rect -51 -64130 996 -64113
rect -67 -64138 -34 -64105
rect -51 -64201 996 -64184
rect -67 -64209 -34 -64176
rect -51 -64272 996 -64255
rect -67 -64280 -34 -64247
rect -51 -64343 996 -64326
rect -67 -64351 -34 -64318
rect -51 -64414 996 -64397
rect -67 -64422 -34 -64389
rect -51 -64485 996 -64468
rect -67 -64493 -34 -64460
rect -51 -64556 996 -64539
rect -67 -64564 -34 -64531
rect -51 -64627 996 -64610
rect -67 -64635 -34 -64602
rect -51 -64698 996 -64681
rect -67 -64706 -34 -64673
rect -51 -64769 996 -64752
rect -67 -64777 -34 -64744
rect -51 -64840 996 -64823
rect -67 -64848 -34 -64815
rect -51 -64911 996 -64894
rect -67 -64919 -34 -64886
rect -51 -64982 996 -64965
rect -67 -64990 -34 -64957
rect -51 -65053 996 -65036
rect -67 -65061 -34 -65028
rect -51 -65124 996 -65107
rect -67 -65132 -34 -65099
rect -51 -65195 996 -65178
rect -67 -65203 -34 -65170
rect -51 -65266 996 -65249
rect -67 -65274 -34 -65241
rect -51 -65337 996 -65320
rect -67 -65345 -34 -65312
rect -51 -65408 996 -65391
rect -67 -65416 -34 -65383
rect -51 -65479 996 -65462
rect -67 -65487 -34 -65454
rect -51 -65550 996 -65533
rect -67 -65558 -34 -65525
rect -51 -65621 996 -65604
rect -67 -65629 -34 -65596
rect -51 -65692 996 -65675
rect -67 -65700 -34 -65667
rect -51 -65763 996 -65746
rect -67 -65771 -34 -65738
rect -51 -65834 996 -65817
rect -67 -65842 -34 -65809
rect -51 -65905 996 -65888
rect -67 -65913 -34 -65880
rect -51 -65976 996 -65959
rect -67 -65984 -34 -65951
rect -51 -66047 996 -66030
rect -67 -66055 -34 -66022
rect -51 -66118 996 -66101
rect -67 -66126 -34 -66093
rect -51 -66189 996 -66172
rect -67 -66197 -34 -66164
rect -51 -66260 996 -66243
rect -67 -66268 -34 -66235
rect -51 -66331 996 -66314
rect -67 -66339 -34 -66306
rect -51 -66402 996 -66385
rect -67 -66410 -34 -66377
rect -51 -66473 996 -66456
rect -67 -66481 -34 -66448
rect -51 -66544 996 -66527
rect -67 -66552 -34 -66519
rect -51 -66615 996 -66598
rect -67 -66623 -34 -66590
rect -51 -66686 996 -66669
rect -67 -66694 -34 -66661
rect -51 -66757 996 -66740
rect -67 -66765 -34 -66732
rect -51 -66828 996 -66811
rect -67 -66836 -34 -66803
rect -51 -66899 996 -66882
rect -67 -66907 -34 -66874
rect -51 -66970 996 -66953
rect -67 -66978 -34 -66945
rect -51 -67041 996 -67024
rect -67 -67049 -34 -67016
rect -51 -67112 996 -67095
rect -67 -67120 -34 -67087
rect -51 -67183 996 -67166
rect -67 -67191 -34 -67158
rect -51 -67254 996 -67237
rect -67 -67262 -34 -67229
rect -51 -67325 996 -67308
rect -67 -67333 -34 -67300
rect -51 -67396 996 -67379
rect -67 -67404 -34 -67371
rect -51 -67467 996 -67450
rect -67 -67475 -34 -67442
rect -51 -67538 996 -67521
rect -67 -67546 -34 -67513
rect -51 -67609 996 -67592
rect -67 -67617 -34 -67584
rect -51 -67680 996 -67663
rect -67 -67688 -34 -67655
rect -51 -67751 996 -67734
rect -67 -67759 -34 -67726
rect -51 -67822 996 -67805
rect -67 -67830 -34 -67797
rect -51 -67893 996 -67876
rect -67 -67901 -34 -67868
rect -51 -67964 996 -67947
rect -67 -67972 -34 -67939
rect -51 -68035 996 -68018
rect -67 -68043 -34 -68010
rect -51 -68106 996 -68089
rect -67 -68114 -34 -68081
rect -51 -68177 996 -68160
rect -67 -68185 -34 -68152
rect -51 -68248 996 -68231
rect -67 -68256 -34 -68223
rect -51 -68319 996 -68302
rect -67 -68327 -34 -68294
rect -51 -68390 996 -68373
rect -67 -68398 -34 -68365
rect -51 -68461 996 -68444
rect -67 -68469 -34 -68436
rect -51 -68532 996 -68515
rect -67 -68540 -34 -68507
rect -51 -68603 996 -68586
rect -67 -68611 -34 -68578
rect -51 -68674 996 -68657
rect -67 -68682 -34 -68649
rect -51 -68745 996 -68728
rect -67 -68753 -34 -68720
rect -51 -68816 996 -68799
rect -67 -68824 -34 -68791
rect -51 -68887 996 -68870
rect -67 -68895 -34 -68862
rect -51 -68958 996 -68941
rect -67 -68966 -34 -68933
rect -51 -69029 996 -69012
rect -67 -69037 -34 -69004
rect -51 -69100 996 -69083
rect -67 -69108 -34 -69075
rect -51 -69171 996 -69154
rect -67 -69179 -34 -69146
rect -51 -69242 996 -69225
rect -67 -69250 -34 -69217
rect -51 -69313 996 -69296
rect -67 -69321 -34 -69288
rect -51 -69384 996 -69367
rect -67 -69392 -34 -69359
rect -51 -69455 996 -69438
rect -67 -69463 -34 -69430
rect -51 -69526 996 -69509
rect -67 -69534 -34 -69501
rect -51 -69597 996 -69580
rect -67 -69605 -34 -69572
rect -51 -69668 996 -69651
rect -67 -69676 -34 -69643
rect -51 -69739 996 -69722
rect -67 -69747 -34 -69714
rect -51 -69810 996 -69793
rect -67 -69818 -34 -69785
rect -51 -69881 996 -69864
rect -67 -69889 -34 -69856
rect -51 -69952 996 -69935
rect -67 -69960 -34 -69927
rect -51 -70023 996 -70006
rect -67 -70031 -34 -69998
rect -51 -70094 996 -70077
rect -67 -70102 -34 -70069
rect -51 -70165 996 -70148
rect -67 -70173 -34 -70140
rect -51 -70236 996 -70219
rect -67 -70244 -34 -70211
rect -51 -70307 996 -70290
rect -67 -70315 -34 -70282
rect -51 -70378 996 -70361
rect -67 -70386 -34 -70353
rect -51 -70449 996 -70432
rect -67 -70457 -34 -70424
rect -51 -70520 996 -70503
rect -67 -70528 -34 -70495
rect -51 -70591 996 -70574
rect -67 -70599 -34 -70566
rect -51 -70662 996 -70645
rect -67 -70670 -34 -70637
rect -51 -70733 996 -70716
rect -67 -70741 -34 -70708
rect -51 -70804 996 -70787
rect -67 -70812 -34 -70779
rect -51 -70875 996 -70858
rect -67 -70883 -34 -70850
rect -51 -70946 996 -70929
rect -67 -70954 -34 -70921
rect -51 -71017 996 -71000
rect -67 -71025 -34 -70992
rect -51 -71088 996 -71071
rect -67 -71096 -34 -71063
rect -51 -71159 996 -71142
rect -67 -71167 -34 -71134
rect -51 -71230 996 -71213
rect -67 -71238 -34 -71205
rect -51 -71301 996 -71284
rect -67 -71309 -34 -71276
rect -51 -71372 996 -71355
rect -67 -71380 -34 -71347
rect -51 -71443 996 -71426
rect -67 -71451 -34 -71418
rect -51 -71514 996 -71497
rect -67 -71522 -34 -71489
rect -51 -71585 996 -71568
rect -67 -71593 -34 -71560
rect -51 -71656 996 -71639
rect -67 -71664 -34 -71631
rect -51 -71727 996 -71710
rect -67 -71735 -34 -71702
rect -51 -71798 996 -71781
rect -67 -71806 -34 -71773
rect -51 -71869 996 -71852
rect -67 -71877 -34 -71844
rect -51 -71940 996 -71923
rect -67 -71948 -34 -71915
rect -51 -72011 996 -71994
rect -67 -72019 -34 -71986
rect -51 -72082 996 -72065
rect -67 -72090 -34 -72057
rect -51 -72153 996 -72136
rect -67 -72161 -34 -72128
rect -51 -72224 996 -72207
rect -67 -72232 -34 -72199
rect -51 -72295 996 -72278
rect -67 -72303 -34 -72270
rect -51 -72366 996 -72349
rect -67 -72374 -34 -72341
rect -51 -72437 996 -72420
rect -67 -72445 -34 -72412
rect -51 -72508 996 -72491
rect -67 -72516 -34 -72483
rect -51 -72579 996 -72562
rect -67 -72587 -34 -72554
rect -51 -72650 996 -72633
rect -67 -72658 -34 -72625
rect -60 166 -27 199
rect -27 174 986 191
<< polycont >>
rect -59 -17 -42 0
rect -59 -88 -42 -71
rect -59 -159 -42 -142
rect -59 -230 -42 -213
rect -59 -301 -42 -284
rect -59 -372 -42 -355
rect -59 -443 -42 -426
rect -59 -514 -42 -497
rect -59 -585 -42 -568
rect -59 -656 -42 -639
rect -59 -727 -42 -710
rect -59 -798 -42 -781
rect -59 -869 -42 -852
rect -59 -940 -42 -923
rect -59 -1011 -42 -994
rect -59 -1082 -42 -1065
rect -59 -1153 -42 -1136
rect -59 -1224 -42 -1207
rect -59 -1295 -42 -1278
rect -59 -1366 -42 -1349
rect -59 -1437 -42 -1420
rect -59 -1508 -42 -1491
rect -59 -1579 -42 -1562
rect -59 -1650 -42 -1633
rect -59 -1721 -42 -1704
rect -59 -1792 -42 -1775
rect -59 -1863 -42 -1846
rect -59 -1934 -42 -1917
rect -59 -2005 -42 -1988
rect -59 -2076 -42 -2059
rect -59 -2147 -42 -2130
rect -59 -2218 -42 -2201
rect -59 -2289 -42 -2272
rect -59 -2360 -42 -2343
rect -59 -2431 -42 -2414
rect -59 -2502 -42 -2485
rect -59 -2573 -42 -2556
rect -59 -2644 -42 -2627
rect -59 -2715 -42 -2698
rect -59 -2786 -42 -2769
rect -59 -2857 -42 -2840
rect -59 -2928 -42 -2911
rect -59 -2999 -42 -2982
rect -59 -3070 -42 -3053
rect -59 -3141 -42 -3124
rect -59 -3212 -42 -3195
rect -59 -3283 -42 -3266
rect -59 -3354 -42 -3337
rect -59 -3425 -42 -3408
rect -59 -3496 -42 -3479
rect -59 -3567 -42 -3550
rect -59 -3638 -42 -3621
rect -59 -3709 -42 -3692
rect -59 -3780 -42 -3763
rect -59 -3851 -42 -3834
rect -59 -3922 -42 -3905
rect -59 -3993 -42 -3976
rect -59 -4064 -42 -4047
rect -59 -4135 -42 -4118
rect -59 -4206 -42 -4189
rect -59 -4277 -42 -4260
rect -59 -4348 -42 -4331
rect -59 -4419 -42 -4402
rect -59 -4490 -42 -4473
rect -59 -4561 -42 -4544
rect -59 -4632 -42 -4615
rect -59 -4703 -42 -4686
rect -59 -4774 -42 -4757
rect -59 -4845 -42 -4828
rect -59 -4916 -42 -4899
rect -59 -4987 -42 -4970
rect -59 -5058 -42 -5041
rect -59 -5129 -42 -5112
rect -59 -5200 -42 -5183
rect -59 -5271 -42 -5254
rect -59 -5342 -42 -5325
rect -59 -5413 -42 -5396
rect -59 -5484 -42 -5467
rect -59 -5555 -42 -5538
rect -59 -5626 -42 -5609
rect -59 -5697 -42 -5680
rect -59 -5768 -42 -5751
rect -59 -5839 -42 -5822
rect -59 -5910 -42 -5893
rect -59 -5981 -42 -5964
rect -59 -6052 -42 -6035
rect -59 -6123 -42 -6106
rect -59 -6194 -42 -6177
rect -59 -6265 -42 -6248
rect -59 -6336 -42 -6319
rect -59 -6407 -42 -6390
rect -59 -6478 -42 -6461
rect -59 -6549 -42 -6532
rect -59 -6620 -42 -6603
rect -59 -6691 -42 -6674
rect -59 -6762 -42 -6745
rect -59 -6833 -42 -6816
rect -59 -6904 -42 -6887
rect -59 -6975 -42 -6958
rect -59 -7046 -42 -7029
rect -59 -7117 -42 -7100
rect -59 -7188 -42 -7171
rect -59 -7259 -42 -7242
rect -59 -7330 -42 -7313
rect -59 -7401 -42 -7384
rect -59 -7472 -42 -7455
rect -59 -7543 -42 -7526
rect -59 -7614 -42 -7597
rect -59 -7685 -42 -7668
rect -59 -7756 -42 -7739
rect -59 -7827 -42 -7810
rect -59 -7898 -42 -7881
rect -59 -7969 -42 -7952
rect -59 -8040 -42 -8023
rect -59 -8111 -42 -8094
rect -59 -8182 -42 -8165
rect -59 -8253 -42 -8236
rect -59 -8324 -42 -8307
rect -59 -8395 -42 -8378
rect -59 -8466 -42 -8449
rect -59 -8537 -42 -8520
rect -59 -8608 -42 -8591
rect -59 -8679 -42 -8662
rect -59 -8750 -42 -8733
rect -59 -8821 -42 -8804
rect -59 -8892 -42 -8875
rect -59 -8963 -42 -8946
rect -59 -9034 -42 -9017
rect -59 -9105 -42 -9088
rect -59 -9176 -42 -9159
rect -59 -9247 -42 -9230
rect -59 -9318 -42 -9301
rect -59 -9389 -42 -9372
rect -59 -9460 -42 -9443
rect -59 -9531 -42 -9514
rect -59 -9602 -42 -9585
rect -59 -9673 -42 -9656
rect -59 -9744 -42 -9727
rect -59 -9815 -42 -9798
rect -59 -9886 -42 -9869
rect -59 -9957 -42 -9940
rect -59 -10028 -42 -10011
rect -59 -10099 -42 -10082
rect -59 -10170 -42 -10153
rect -59 -10241 -42 -10224
rect -59 -10312 -42 -10295
rect -59 -10383 -42 -10366
rect -59 -10454 -42 -10437
rect -59 -10525 -42 -10508
rect -59 -10596 -42 -10579
rect -59 -10667 -42 -10650
rect -59 -10738 -42 -10721
rect -59 -10809 -42 -10792
rect -59 -10880 -42 -10863
rect -59 -10951 -42 -10934
rect -59 -11022 -42 -11005
rect -59 -11093 -42 -11076
rect -59 -11164 -42 -11147
rect -59 -11235 -42 -11218
rect -59 -11306 -42 -11289
rect -59 -11377 -42 -11360
rect -59 -11448 -42 -11431
rect -59 -11519 -42 -11502
rect -59 -11590 -42 -11573
rect -59 -11661 -42 -11644
rect -59 -11732 -42 -11715
rect -59 -11803 -42 -11786
rect -59 -11874 -42 -11857
rect -59 -11945 -42 -11928
rect -59 -12016 -42 -11999
rect -59 -12087 -42 -12070
rect -59 -12158 -42 -12141
rect -59 -12229 -42 -12212
rect -59 -12300 -42 -12283
rect -59 -12371 -42 -12354
rect -59 -12442 -42 -12425
rect -59 -12513 -42 -12496
rect -59 -12584 -42 -12567
rect -59 -12655 -42 -12638
rect -59 -12726 -42 -12709
rect -59 -12797 -42 -12780
rect -59 -12868 -42 -12851
rect -59 -12939 -42 -12922
rect -59 -13010 -42 -12993
rect -59 -13081 -42 -13064
rect -59 -13152 -42 -13135
rect -59 -13223 -42 -13206
rect -59 -13294 -42 -13277
rect -59 -13365 -42 -13348
rect -59 -13436 -42 -13419
rect -59 -13507 -42 -13490
rect -59 -13578 -42 -13561
rect -59 -13649 -42 -13632
rect -59 -13720 -42 -13703
rect -59 -13791 -42 -13774
rect -59 -13862 -42 -13845
rect -59 -13933 -42 -13916
rect -59 -14004 -42 -13987
rect -59 -14075 -42 -14058
rect -59 -14146 -42 -14129
rect -59 -14217 -42 -14200
rect -59 -14288 -42 -14271
rect -59 -14359 -42 -14342
rect -59 -14430 -42 -14413
rect -59 -14501 -42 -14484
rect -59 -14572 -42 -14555
rect -59 -14643 -42 -14626
rect -59 -14714 -42 -14697
rect -59 -14785 -42 -14768
rect -59 -14856 -42 -14839
rect -59 -14927 -42 -14910
rect -59 -14998 -42 -14981
rect -59 -15069 -42 -15052
rect -59 -15140 -42 -15123
rect -59 -15211 -42 -15194
rect -59 -15282 -42 -15265
rect -59 -15353 -42 -15336
rect -59 -15424 -42 -15407
rect -59 -15495 -42 -15478
rect -59 -15566 -42 -15549
rect -59 -15637 -42 -15620
rect -59 -15708 -42 -15691
rect -59 -15779 -42 -15762
rect -59 -15850 -42 -15833
rect -59 -15921 -42 -15904
rect -59 -15992 -42 -15975
rect -59 -16063 -42 -16046
rect -59 -16134 -42 -16117
rect -59 -16205 -42 -16188
rect -59 -16276 -42 -16259
rect -59 -16347 -42 -16330
rect -59 -16418 -42 -16401
rect -59 -16489 -42 -16472
rect -59 -16560 -42 -16543
rect -59 -16631 -42 -16614
rect -59 -16702 -42 -16685
rect -59 -16773 -42 -16756
rect -59 -16844 -42 -16827
rect -59 -16915 -42 -16898
rect -59 -16986 -42 -16969
rect -59 -17057 -42 -17040
rect -59 -17128 -42 -17111
rect -59 -17199 -42 -17182
rect -59 -17270 -42 -17253
rect -59 -17341 -42 -17324
rect -59 -17412 -42 -17395
rect -59 -17483 -42 -17466
rect -59 -17554 -42 -17537
rect -59 -17625 -42 -17608
rect -59 -17696 -42 -17679
rect -59 -17767 -42 -17750
rect -59 -17838 -42 -17821
rect -59 -17909 -42 -17892
rect -59 -17980 -42 -17963
rect -59 -18051 -42 -18034
rect -59 -18122 -42 -18105
rect -59 -18193 -42 -18176
rect -59 -18264 -42 -18247
rect -59 -18335 -42 -18318
rect -59 -18406 -42 -18389
rect -59 -18477 -42 -18460
rect -59 -18548 -42 -18531
rect -59 -18619 -42 -18602
rect -59 -18690 -42 -18673
rect -59 -18761 -42 -18744
rect -59 -18832 -42 -18815
rect -59 -18903 -42 -18886
rect -59 -18974 -42 -18957
rect -59 -19045 -42 -19028
rect -59 -19116 -42 -19099
rect -59 -19187 -42 -19170
rect -59 -19258 -42 -19241
rect -59 -19329 -42 -19312
rect -59 -19400 -42 -19383
rect -59 -19471 -42 -19454
rect -59 -19542 -42 -19525
rect -59 -19613 -42 -19596
rect -59 -19684 -42 -19667
rect -59 -19755 -42 -19738
rect -59 -19826 -42 -19809
rect -59 -19897 -42 -19880
rect -59 -19968 -42 -19951
rect -59 -20039 -42 -20022
rect -59 -20110 -42 -20093
rect -59 -20181 -42 -20164
rect -59 -20252 -42 -20235
rect -59 -20323 -42 -20306
rect -59 -20394 -42 -20377
rect -59 -20465 -42 -20448
rect -59 -20536 -42 -20519
rect -59 -20607 -42 -20590
rect -59 -20678 -42 -20661
rect -59 -20749 -42 -20732
rect -59 -20820 -42 -20803
rect -59 -20891 -42 -20874
rect -59 -20962 -42 -20945
rect -59 -21033 -42 -21016
rect -59 -21104 -42 -21087
rect -59 -21175 -42 -21158
rect -59 -21246 -42 -21229
rect -59 -21317 -42 -21300
rect -59 -21388 -42 -21371
rect -59 -21459 -42 -21442
rect -59 -21530 -42 -21513
rect -59 -21601 -42 -21584
rect -59 -21672 -42 -21655
rect -59 -21743 -42 -21726
rect -59 -21814 -42 -21797
rect -59 -21885 -42 -21868
rect -59 -21956 -42 -21939
rect -59 -22027 -42 -22010
rect -59 -22098 -42 -22081
rect -59 -22169 -42 -22152
rect -59 -22240 -42 -22223
rect -59 -22311 -42 -22294
rect -59 -22382 -42 -22365
rect -59 -22453 -42 -22436
rect -59 -22524 -42 -22507
rect -59 -22595 -42 -22578
rect -59 -22666 -42 -22649
rect -59 -22737 -42 -22720
rect -59 -22808 -42 -22791
rect -59 -22879 -42 -22862
rect -59 -22950 -42 -22933
rect -59 -23021 -42 -23004
rect -59 -23092 -42 -23075
rect -59 -23163 -42 -23146
rect -59 -23234 -42 -23217
rect -59 -23305 -42 -23288
rect -59 -23376 -42 -23359
rect -59 -23447 -42 -23430
rect -59 -23518 -42 -23501
rect -59 -23589 -42 -23572
rect -59 -23660 -42 -23643
rect -59 -23731 -42 -23714
rect -59 -23802 -42 -23785
rect -59 -23873 -42 -23856
rect -59 -23944 -42 -23927
rect -59 -24015 -42 -23998
rect -59 -24086 -42 -24069
rect -59 -24157 -42 -24140
rect -59 -24228 -42 -24211
rect -59 -24299 -42 -24282
rect -59 -24370 -42 -24353
rect -59 -24441 -42 -24424
rect -59 -24512 -42 -24495
rect -59 -24583 -42 -24566
rect -59 -24654 -42 -24637
rect -59 -24725 -42 -24708
rect -59 -24796 -42 -24779
rect -59 -24867 -42 -24850
rect -59 -24938 -42 -24921
rect -59 -25009 -42 -24992
rect -59 -25080 -42 -25063
rect -59 -25151 -42 -25134
rect -59 -25222 -42 -25205
rect -59 -25293 -42 -25276
rect -59 -25364 -42 -25347
rect -59 -25435 -42 -25418
rect -59 -25506 -42 -25489
rect -59 -25577 -42 -25560
rect -59 -25648 -42 -25631
rect -59 -25719 -42 -25702
rect -59 -25790 -42 -25773
rect -59 -25861 -42 -25844
rect -59 -25932 -42 -25915
rect -59 -26003 -42 -25986
rect -59 -26074 -42 -26057
rect -59 -26145 -42 -26128
rect -59 -26216 -42 -26199
rect -59 -26287 -42 -26270
rect -59 -26358 -42 -26341
rect -59 -26429 -42 -26412
rect -59 -26500 -42 -26483
rect -59 -26571 -42 -26554
rect -59 -26642 -42 -26625
rect -59 -26713 -42 -26696
rect -59 -26784 -42 -26767
rect -59 -26855 -42 -26838
rect -59 -26926 -42 -26909
rect -59 -26997 -42 -26980
rect -59 -27068 -42 -27051
rect -59 -27139 -42 -27122
rect -59 -27210 -42 -27193
rect -59 -27281 -42 -27264
rect -59 -27352 -42 -27335
rect -59 -27423 -42 -27406
rect -59 -27494 -42 -27477
rect -59 -27565 -42 -27548
rect -59 -27636 -42 -27619
rect -59 -27707 -42 -27690
rect -59 -27778 -42 -27761
rect -59 -27849 -42 -27832
rect -59 -27920 -42 -27903
rect -59 -27991 -42 -27974
rect -59 -28062 -42 -28045
rect -59 -28133 -42 -28116
rect -59 -28204 -42 -28187
rect -59 -28275 -42 -28258
rect -59 -28346 -42 -28329
rect -59 -28417 -42 -28400
rect -59 -28488 -42 -28471
rect -59 -28559 -42 -28542
rect -59 -28630 -42 -28613
rect -59 -28701 -42 -28684
rect -59 -28772 -42 -28755
rect -59 -28843 -42 -28826
rect -59 -28914 -42 -28897
rect -59 -28985 -42 -28968
rect -59 -29056 -42 -29039
rect -59 -29127 -42 -29110
rect -59 -29198 -42 -29181
rect -59 -29269 -42 -29252
rect -59 -29340 -42 -29323
rect -59 -29411 -42 -29394
rect -59 -29482 -42 -29465
rect -59 -29553 -42 -29536
rect -59 -29624 -42 -29607
rect -59 -29695 -42 -29678
rect -59 -29766 -42 -29749
rect -59 -29837 -42 -29820
rect -59 -29908 -42 -29891
rect -59 -29979 -42 -29962
rect -59 -30050 -42 -30033
rect -59 -30121 -42 -30104
rect -59 -30192 -42 -30175
rect -59 -30263 -42 -30246
rect -59 -30334 -42 -30317
rect -59 -30405 -42 -30388
rect -59 -30476 -42 -30459
rect -59 -30547 -42 -30530
rect -59 -30618 -42 -30601
rect -59 -30689 -42 -30672
rect -59 -30760 -42 -30743
rect -59 -30831 -42 -30814
rect -59 -30902 -42 -30885
rect -59 -30973 -42 -30956
rect -59 -31044 -42 -31027
rect -59 -31115 -42 -31098
rect -59 -31186 -42 -31169
rect -59 -31257 -42 -31240
rect -59 -31328 -42 -31311
rect -59 -31399 -42 -31382
rect -59 -31470 -42 -31453
rect -59 -31541 -42 -31524
rect -59 -31612 -42 -31595
rect -59 -31683 -42 -31666
rect -59 -31754 -42 -31737
rect -59 -31825 -42 -31808
rect -59 -31896 -42 -31879
rect -59 -31967 -42 -31950
rect -59 -32038 -42 -32021
rect -59 -32109 -42 -32092
rect -59 -32180 -42 -32163
rect -59 -32251 -42 -32234
rect -59 -32322 -42 -32305
rect -59 -32393 -42 -32376
rect -59 -32464 -42 -32447
rect -59 -32535 -42 -32518
rect -59 -32606 -42 -32589
rect -59 -32677 -42 -32660
rect -59 -32748 -42 -32731
rect -59 -32819 -42 -32802
rect -59 -32890 -42 -32873
rect -59 -32961 -42 -32944
rect -59 -33032 -42 -33015
rect -59 -33103 -42 -33086
rect -59 -33174 -42 -33157
rect -59 -33245 -42 -33228
rect -59 -33316 -42 -33299
rect -59 -33387 -42 -33370
rect -59 -33458 -42 -33441
rect -59 -33529 -42 -33512
rect -59 -33600 -42 -33583
rect -59 -33671 -42 -33654
rect -59 -33742 -42 -33725
rect -59 -33813 -42 -33796
rect -59 -33884 -42 -33867
rect -59 -33955 -42 -33938
rect -59 -34026 -42 -34009
rect -59 -34097 -42 -34080
rect -59 -34168 -42 -34151
rect -59 -34239 -42 -34222
rect -59 -34310 -42 -34293
rect -59 -34381 -42 -34364
rect -59 -34452 -42 -34435
rect -59 -34523 -42 -34506
rect -59 -34594 -42 -34577
rect -59 -34665 -42 -34648
rect -59 -34736 -42 -34719
rect -59 -34807 -42 -34790
rect -59 -34878 -42 -34861
rect -59 -34949 -42 -34932
rect -59 -35020 -42 -35003
rect -59 -35091 -42 -35074
rect -59 -35162 -42 -35145
rect -59 -35233 -42 -35216
rect -59 -35304 -42 -35287
rect -59 -35375 -42 -35358
rect -59 -35446 -42 -35429
rect -59 -35517 -42 -35500
rect -59 -35588 -42 -35571
rect -59 -35659 -42 -35642
rect -59 -35730 -42 -35713
rect -59 -35801 -42 -35784
rect -59 -35872 -42 -35855
rect -59 -35943 -42 -35926
rect -59 -36014 -42 -35997
rect -59 -36085 -42 -36068
rect -59 -36156 -42 -36139
rect -59 -36227 -42 -36210
rect -59 -36298 -42 -36281
rect -59 -36369 -42 -36352
rect -59 -36440 -42 -36423
rect -59 -36511 -42 -36494
rect -59 -36582 -42 -36565
rect -59 -36653 -42 -36636
rect -59 -36724 -42 -36707
rect -59 -36795 -42 -36778
rect -59 -36866 -42 -36849
rect -59 -36937 -42 -36920
rect -59 -37008 -42 -36991
rect -59 -37079 -42 -37062
rect -59 -37150 -42 -37133
rect -59 -37221 -42 -37204
rect -59 -37292 -42 -37275
rect -59 -37363 -42 -37346
rect -59 -37434 -42 -37417
rect -59 -37505 -42 -37488
rect -59 -37576 -42 -37559
rect -59 -37647 -42 -37630
rect -59 -37718 -42 -37701
rect -59 -37789 -42 -37772
rect -59 -37860 -42 -37843
rect -59 -37931 -42 -37914
rect -59 -38002 -42 -37985
rect -59 -38073 -42 -38056
rect -59 -38144 -42 -38127
rect -59 -38215 -42 -38198
rect -59 -38286 -42 -38269
rect -59 -38357 -42 -38340
rect -59 -38428 -42 -38411
rect -59 -38499 -42 -38482
rect -59 -38570 -42 -38553
rect -59 -38641 -42 -38624
rect -59 -38712 -42 -38695
rect -59 -38783 -42 -38766
rect -59 -38854 -42 -38837
rect -59 -38925 -42 -38908
rect -59 -38996 -42 -38979
rect -59 -39067 -42 -39050
rect -59 -39138 -42 -39121
rect -59 -39209 -42 -39192
rect -59 -39280 -42 -39263
rect -59 -39351 -42 -39334
rect -59 -39422 -42 -39405
rect -59 -39493 -42 -39476
rect -59 -39564 -42 -39547
rect -59 -39635 -42 -39618
rect -59 -39706 -42 -39689
rect -59 -39777 -42 -39760
rect -59 -39848 -42 -39831
rect -59 -39919 -42 -39902
rect -59 -39990 -42 -39973
rect -59 -40061 -42 -40044
rect -59 -40132 -42 -40115
rect -59 -40203 -42 -40186
rect -59 -40274 -42 -40257
rect -59 -40345 -42 -40328
rect -59 -40416 -42 -40399
rect -59 -40487 -42 -40470
rect -59 -40558 -42 -40541
rect -59 -40629 -42 -40612
rect -59 -40700 -42 -40683
rect -59 -40771 -42 -40754
rect -59 -40842 -42 -40825
rect -59 -40913 -42 -40896
rect -59 -40984 -42 -40967
rect -59 -41055 -42 -41038
rect -59 -41126 -42 -41109
rect -59 -41197 -42 -41180
rect -59 -41268 -42 -41251
rect -59 -41339 -42 -41322
rect -59 -41410 -42 -41393
rect -59 -41481 -42 -41464
rect -59 -41552 -42 -41535
rect -59 -41623 -42 -41606
rect -59 -41694 -42 -41677
rect -59 -41765 -42 -41748
rect -59 -41836 -42 -41819
rect -59 -41907 -42 -41890
rect -59 -41978 -42 -41961
rect -59 -42049 -42 -42032
rect -59 -42120 -42 -42103
rect -59 -42191 -42 -42174
rect -59 -42262 -42 -42245
rect -59 -42333 -42 -42316
rect -59 -42404 -42 -42387
rect -59 -42475 -42 -42458
rect -59 -42546 -42 -42529
rect -59 -42617 -42 -42600
rect -59 -42688 -42 -42671
rect -59 -42759 -42 -42742
rect -59 -42830 -42 -42813
rect -59 -42901 -42 -42884
rect -59 -42972 -42 -42955
rect -59 -43043 -42 -43026
rect -59 -43114 -42 -43097
rect -59 -43185 -42 -43168
rect -59 -43256 -42 -43239
rect -59 -43327 -42 -43310
rect -59 -43398 -42 -43381
rect -59 -43469 -42 -43452
rect -59 -43540 -42 -43523
rect -59 -43611 -42 -43594
rect -59 -43682 -42 -43665
rect -59 -43753 -42 -43736
rect -59 -43824 -42 -43807
rect -59 -43895 -42 -43878
rect -59 -43966 -42 -43949
rect -59 -44037 -42 -44020
rect -59 -44108 -42 -44091
rect -59 -44179 -42 -44162
rect -59 -44250 -42 -44233
rect -59 -44321 -42 -44304
rect -59 -44392 -42 -44375
rect -59 -44463 -42 -44446
rect -59 -44534 -42 -44517
rect -59 -44605 -42 -44588
rect -59 -44676 -42 -44659
rect -59 -44747 -42 -44730
rect -59 -44818 -42 -44801
rect -59 -44889 -42 -44872
rect -59 -44960 -42 -44943
rect -59 -45031 -42 -45014
rect -59 -45102 -42 -45085
rect -59 -45173 -42 -45156
rect -59 -45244 -42 -45227
rect -59 -45315 -42 -45298
rect -59 -45386 -42 -45369
rect -59 -45457 -42 -45440
rect -59 -45528 -42 -45511
rect -59 -45599 -42 -45582
rect -59 -45670 -42 -45653
rect -59 -45741 -42 -45724
rect -59 -45812 -42 -45795
rect -59 -45883 -42 -45866
rect -59 -45954 -42 -45937
rect -59 -46025 -42 -46008
rect -59 -46096 -42 -46079
rect -59 -46167 -42 -46150
rect -59 -46238 -42 -46221
rect -59 -46309 -42 -46292
rect -59 -46380 -42 -46363
rect -59 -46451 -42 -46434
rect -59 -46522 -42 -46505
rect -59 -46593 -42 -46576
rect -59 -46664 -42 -46647
rect -59 -46735 -42 -46718
rect -59 -46806 -42 -46789
rect -59 -46877 -42 -46860
rect -59 -46948 -42 -46931
rect -59 -47019 -42 -47002
rect -59 -47090 -42 -47073
rect -59 -47161 -42 -47144
rect -59 -47232 -42 -47215
rect -59 -47303 -42 -47286
rect -59 -47374 -42 -47357
rect -59 -47445 -42 -47428
rect -59 -47516 -42 -47499
rect -59 -47587 -42 -47570
rect -59 -47658 -42 -47641
rect -59 -47729 -42 -47712
rect -59 -47800 -42 -47783
rect -59 -47871 -42 -47854
rect -59 -47942 -42 -47925
rect -59 -48013 -42 -47996
rect -59 -48084 -42 -48067
rect -59 -48155 -42 -48138
rect -59 -48226 -42 -48209
rect -59 -48297 -42 -48280
rect -59 -48368 -42 -48351
rect -59 -48439 -42 -48422
rect -59 -48510 -42 -48493
rect -59 -48581 -42 -48564
rect -59 -48652 -42 -48635
rect -59 -48723 -42 -48706
rect -59 -48794 -42 -48777
rect -59 -48865 -42 -48848
rect -59 -48936 -42 -48919
rect -59 -49007 -42 -48990
rect -59 -49078 -42 -49061
rect -59 -49149 -42 -49132
rect -59 -49220 -42 -49203
rect -59 -49291 -42 -49274
rect -59 -49362 -42 -49345
rect -59 -49433 -42 -49416
rect -59 -49504 -42 -49487
rect -59 -49575 -42 -49558
rect -59 -49646 -42 -49629
rect -59 -49717 -42 -49700
rect -59 -49788 -42 -49771
rect -59 -49859 -42 -49842
rect -59 -49930 -42 -49913
rect -59 -50001 -42 -49984
rect -59 -50072 -42 -50055
rect -59 -50143 -42 -50126
rect -59 -50214 -42 -50197
rect -59 -50285 -42 -50268
rect -59 -50356 -42 -50339
rect -59 -50427 -42 -50410
rect -59 -50498 -42 -50481
rect -59 -50569 -42 -50552
rect -59 -50640 -42 -50623
rect -59 -50711 -42 -50694
rect -59 -50782 -42 -50765
rect -59 -50853 -42 -50836
rect -59 -50924 -42 -50907
rect -59 -50995 -42 -50978
rect -59 -51066 -42 -51049
rect -59 -51137 -42 -51120
rect -59 -51208 -42 -51191
rect -59 -51279 -42 -51262
rect -59 -51350 -42 -51333
rect -59 -51421 -42 -51404
rect -59 -51492 -42 -51475
rect -59 -51563 -42 -51546
rect -59 -51634 -42 -51617
rect -59 -51705 -42 -51688
rect -59 -51776 -42 -51759
rect -59 -51847 -42 -51830
rect -59 -51918 -42 -51901
rect -59 -51989 -42 -51972
rect -59 -52060 -42 -52043
rect -59 -52131 -42 -52114
rect -59 -52202 -42 -52185
rect -59 -52273 -42 -52256
rect -59 -52344 -42 -52327
rect -59 -52415 -42 -52398
rect -59 -52486 -42 -52469
rect -59 -52557 -42 -52540
rect -59 -52628 -42 -52611
rect -59 -52699 -42 -52682
rect -59 -52770 -42 -52753
rect -59 -52841 -42 -52824
rect -59 -52912 -42 -52895
rect -59 -52983 -42 -52966
rect -59 -53054 -42 -53037
rect -59 -53125 -42 -53108
rect -59 -53196 -42 -53179
rect -59 -53267 -42 -53250
rect -59 -53338 -42 -53321
rect -59 -53409 -42 -53392
rect -59 -53480 -42 -53463
rect -59 -53551 -42 -53534
rect -59 -53622 -42 -53605
rect -59 -53693 -42 -53676
rect -59 -53764 -42 -53747
rect -59 -53835 -42 -53818
rect -59 -53906 -42 -53889
rect -59 -53977 -42 -53960
rect -59 -54048 -42 -54031
rect -59 -54119 -42 -54102
rect -59 -54190 -42 -54173
rect -59 -54261 -42 -54244
rect -59 -54332 -42 -54315
rect -59 -54403 -42 -54386
rect -59 -54474 -42 -54457
rect -59 -54545 -42 -54528
rect -59 -54616 -42 -54599
rect -59 -54687 -42 -54670
rect -59 -54758 -42 -54741
rect -59 -54829 -42 -54812
rect -59 -54900 -42 -54883
rect -59 -54971 -42 -54954
rect -59 -55042 -42 -55025
rect -59 -55113 -42 -55096
rect -59 -55184 -42 -55167
rect -59 -55255 -42 -55238
rect -59 -55326 -42 -55309
rect -59 -55397 -42 -55380
rect -59 -55468 -42 -55451
rect -59 -55539 -42 -55522
rect -59 -55610 -42 -55593
rect -59 -55681 -42 -55664
rect -59 -55752 -42 -55735
rect -59 -55823 -42 -55806
rect -59 -55894 -42 -55877
rect -59 -55965 -42 -55948
rect -59 -56036 -42 -56019
rect -59 -56107 -42 -56090
rect -59 -56178 -42 -56161
rect -59 -56249 -42 -56232
rect -59 -56320 -42 -56303
rect -59 -56391 -42 -56374
rect -59 -56462 -42 -56445
rect -59 -56533 -42 -56516
rect -59 -56604 -42 -56587
rect -59 -56675 -42 -56658
rect -59 -56746 -42 -56729
rect -59 -56817 -42 -56800
rect -59 -56888 -42 -56871
rect -59 -56959 -42 -56942
rect -59 -57030 -42 -57013
rect -59 -57101 -42 -57084
rect -59 -57172 -42 -57155
rect -59 -57243 -42 -57226
rect -59 -57314 -42 -57297
rect -59 -57385 -42 -57368
rect -59 -57456 -42 -57439
rect -59 -57527 -42 -57510
rect -59 -57598 -42 -57581
rect -59 -57669 -42 -57652
rect -59 -57740 -42 -57723
rect -59 -57811 -42 -57794
rect -59 -57882 -42 -57865
rect -59 -57953 -42 -57936
rect -59 -58024 -42 -58007
rect -59 -58095 -42 -58078
rect -59 -58166 -42 -58149
rect -59 -58237 -42 -58220
rect -59 -58308 -42 -58291
rect -59 -58379 -42 -58362
rect -59 -58450 -42 -58433
rect -59 -58521 -42 -58504
rect -59 -58592 -42 -58575
rect -59 -58663 -42 -58646
rect -59 -58734 -42 -58717
rect -59 -58805 -42 -58788
rect -59 -58876 -42 -58859
rect -59 -58947 -42 -58930
rect -59 -59018 -42 -59001
rect -59 -59089 -42 -59072
rect -59 -59160 -42 -59143
rect -59 -59231 -42 -59214
rect -59 -59302 -42 -59285
rect -59 -59373 -42 -59356
rect -59 -59444 -42 -59427
rect -59 -59515 -42 -59498
rect -59 -59586 -42 -59569
rect -59 -59657 -42 -59640
rect -59 -59728 -42 -59711
rect -59 -59799 -42 -59782
rect -59 -59870 -42 -59853
rect -59 -59941 -42 -59924
rect -59 -60012 -42 -59995
rect -59 -60083 -42 -60066
rect -59 -60154 -42 -60137
rect -59 -60225 -42 -60208
rect -59 -60296 -42 -60279
rect -59 -60367 -42 -60350
rect -59 -60438 -42 -60421
rect -59 -60509 -42 -60492
rect -59 -60580 -42 -60563
rect -59 -60651 -42 -60634
rect -59 -60722 -42 -60705
rect -59 -60793 -42 -60776
rect -59 -60864 -42 -60847
rect -59 -60935 -42 -60918
rect -59 -61006 -42 -60989
rect -59 -61077 -42 -61060
rect -59 -61148 -42 -61131
rect -59 -61219 -42 -61202
rect -59 -61290 -42 -61273
rect -59 -61361 -42 -61344
rect -59 -61432 -42 -61415
rect -59 -61503 -42 -61486
rect -59 -61574 -42 -61557
rect -59 -61645 -42 -61628
rect -59 -61716 -42 -61699
rect -59 -61787 -42 -61770
rect -59 -61858 -42 -61841
rect -59 -61929 -42 -61912
rect -59 -62000 -42 -61983
rect -59 -62071 -42 -62054
rect -59 -62142 -42 -62125
rect -59 -62213 -42 -62196
rect -59 -62284 -42 -62267
rect -59 -62355 -42 -62338
rect -59 -62426 -42 -62409
rect -59 -62497 -42 -62480
rect -59 -62568 -42 -62551
rect -59 -62639 -42 -62622
rect -59 -62710 -42 -62693
rect -59 -62781 -42 -62764
rect -59 -62852 -42 -62835
rect -59 -62923 -42 -62906
rect -59 -62994 -42 -62977
rect -59 -63065 -42 -63048
rect -59 -63136 -42 -63119
rect -59 -63207 -42 -63190
rect -59 -63278 -42 -63261
rect -59 -63349 -42 -63332
rect -59 -63420 -42 -63403
rect -59 -63491 -42 -63474
rect -59 -63562 -42 -63545
rect -59 -63633 -42 -63616
rect -59 -63704 -42 -63687
rect -59 -63775 -42 -63758
rect -59 -63846 -42 -63829
rect -59 -63917 -42 -63900
rect -59 -63988 -42 -63971
rect -59 -64059 -42 -64042
rect -59 -64130 -42 -64113
rect -59 -64201 -42 -64184
rect -59 -64272 -42 -64255
rect -59 -64343 -42 -64326
rect -59 -64414 -42 -64397
rect -59 -64485 -42 -64468
rect -59 -64556 -42 -64539
rect -59 -64627 -42 -64610
rect -59 -64698 -42 -64681
rect -59 -64769 -42 -64752
rect -59 -64840 -42 -64823
rect -59 -64911 -42 -64894
rect -59 -64982 -42 -64965
rect -59 -65053 -42 -65036
rect -59 -65124 -42 -65107
rect -59 -65195 -42 -65178
rect -59 -65266 -42 -65249
rect -59 -65337 -42 -65320
rect -59 -65408 -42 -65391
rect -59 -65479 -42 -65462
rect -59 -65550 -42 -65533
rect -59 -65621 -42 -65604
rect -59 -65692 -42 -65675
rect -59 -65763 -42 -65746
rect -59 -65834 -42 -65817
rect -59 -65905 -42 -65888
rect -59 -65976 -42 -65959
rect -59 -66047 -42 -66030
rect -59 -66118 -42 -66101
rect -59 -66189 -42 -66172
rect -59 -66260 -42 -66243
rect -59 -66331 -42 -66314
rect -59 -66402 -42 -66385
rect -59 -66473 -42 -66456
rect -59 -66544 -42 -66527
rect -59 -66615 -42 -66598
rect -59 -66686 -42 -66669
rect -59 -66757 -42 -66740
rect -59 -66828 -42 -66811
rect -59 -66899 -42 -66882
rect -59 -66970 -42 -66953
rect -59 -67041 -42 -67024
rect -59 -67112 -42 -67095
rect -59 -67183 -42 -67166
rect -59 -67254 -42 -67237
rect -59 -67325 -42 -67308
rect -59 -67396 -42 -67379
rect -59 -67467 -42 -67450
rect -59 -67538 -42 -67521
rect -59 -67609 -42 -67592
rect -59 -67680 -42 -67663
rect -59 -67751 -42 -67734
rect -59 -67822 -42 -67805
rect -59 -67893 -42 -67876
rect -59 -67964 -42 -67947
rect -59 -68035 -42 -68018
rect -59 -68106 -42 -68089
rect -59 -68177 -42 -68160
rect -59 -68248 -42 -68231
rect -59 -68319 -42 -68302
rect -59 -68390 -42 -68373
rect -59 -68461 -42 -68444
rect -59 -68532 -42 -68515
rect -59 -68603 -42 -68586
rect -59 -68674 -42 -68657
rect -59 -68745 -42 -68728
rect -59 -68816 -42 -68799
rect -59 -68887 -42 -68870
rect -59 -68958 -42 -68941
rect -59 -69029 -42 -69012
rect -59 -69100 -42 -69083
rect -59 -69171 -42 -69154
rect -59 -69242 -42 -69225
rect -59 -69313 -42 -69296
rect -59 -69384 -42 -69367
rect -59 -69455 -42 -69438
rect -59 -69526 -42 -69509
rect -59 -69597 -42 -69580
rect -59 -69668 -42 -69651
rect -59 -69739 -42 -69722
rect -59 -69810 -42 -69793
rect -59 -69881 -42 -69864
rect -59 -69952 -42 -69935
rect -59 -70023 -42 -70006
rect -59 -70094 -42 -70077
rect -59 -70165 -42 -70148
rect -59 -70236 -42 -70219
rect -59 -70307 -42 -70290
rect -59 -70378 -42 -70361
rect -59 -70449 -42 -70432
rect -59 -70520 -42 -70503
rect -59 -70591 -42 -70574
rect -59 -70662 -42 -70645
rect -59 -70733 -42 -70716
rect -59 -70804 -42 -70787
rect -59 -70875 -42 -70858
rect -59 -70946 -42 -70929
rect -59 -71017 -42 -71000
rect -59 -71088 -42 -71071
rect -59 -71159 -42 -71142
rect -59 -71230 -42 -71213
rect -59 -71301 -42 -71284
rect -59 -71372 -42 -71355
rect -59 -71443 -42 -71426
rect -59 -71514 -42 -71497
rect -59 -71585 -42 -71568
rect -59 -71656 -42 -71639
rect -59 -71727 -42 -71710
rect -59 -71798 -42 -71781
rect -59 -71869 -42 -71852
rect -59 -71940 -42 -71923
rect -59 -72011 -42 -71994
rect -59 -72082 -42 -72065
rect -59 -72153 -42 -72136
rect -59 -72224 -42 -72207
rect -59 -72295 -42 -72278
rect -59 -72366 -42 -72349
rect -59 -72437 -42 -72420
rect -59 -72508 -42 -72491
rect -59 -72579 -42 -72562
rect -59 -72650 -42 -72633
rect -52 174 -35 191
<< locali >>
rect -67 -25 -34 8
rect -67 -96 -34 -63
rect -67 -167 -34 -134
rect -67 -238 -34 -205
rect -67 -309 -34 -276
rect -67 -380 -34 -347
rect -67 -451 -34 -418
rect -67 -522 -34 -489
rect -67 -593 -34 -560
rect -67 -664 -34 -631
rect -67 -735 -34 -702
rect -67 -806 -34 -773
rect -67 -877 -34 -844
rect -67 -948 -34 -915
rect -67 -1019 -34 -986
rect -67 -1090 -34 -1057
rect -67 -1161 -34 -1128
rect -67 -1232 -34 -1199
rect -67 -1303 -34 -1270
rect -67 -1374 -34 -1341
rect -67 -1445 -34 -1412
rect -67 -1516 -34 -1483
rect -67 -1587 -34 -1554
rect -67 -1658 -34 -1625
rect -67 -1729 -34 -1696
rect -67 -1800 -34 -1767
rect -67 -1871 -34 -1838
rect -67 -1942 -34 -1909
rect -67 -2013 -34 -1980
rect -67 -2084 -34 -2051
rect -67 -2155 -34 -2122
rect -67 -2226 -34 -2193
rect -67 -2297 -34 -2264
rect -67 -2368 -34 -2335
rect -67 -2439 -34 -2406
rect -67 -2510 -34 -2477
rect -67 -2581 -34 -2548
rect -67 -2652 -34 -2619
rect -67 -2723 -34 -2690
rect -67 -2794 -34 -2761
rect -67 -2865 -34 -2832
rect -67 -2936 -34 -2903
rect -67 -3007 -34 -2974
rect -67 -3078 -34 -3045
rect -67 -3149 -34 -3116
rect -67 -3220 -34 -3187
rect -67 -3291 -34 -3258
rect -67 -3362 -34 -3329
rect -67 -3433 -34 -3400
rect -67 -3504 -34 -3471
rect -67 -3575 -34 -3542
rect -67 -3646 -34 -3613
rect -67 -3717 -34 -3684
rect -67 -3788 -34 -3755
rect -67 -3859 -34 -3826
rect -67 -3930 -34 -3897
rect -67 -4001 -34 -3968
rect -67 -4072 -34 -4039
rect -67 -4143 -34 -4110
rect -67 -4214 -34 -4181
rect -67 -4285 -34 -4252
rect -67 -4356 -34 -4323
rect -67 -4427 -34 -4394
rect -67 -4498 -34 -4465
rect -67 -4569 -34 -4536
rect -67 -4640 -34 -4607
rect -67 -4711 -34 -4678
rect -67 -4782 -34 -4749
rect -67 -4853 -34 -4820
rect -67 -4924 -34 -4891
rect -67 -4995 -34 -4962
rect -67 -5066 -34 -5033
rect -67 -5137 -34 -5104
rect -67 -5208 -34 -5175
rect -67 -5279 -34 -5246
rect -67 -5350 -34 -5317
rect -67 -5421 -34 -5388
rect -67 -5492 -34 -5459
rect -67 -5563 -34 -5530
rect -67 -5634 -34 -5601
rect -67 -5705 -34 -5672
rect -67 -5776 -34 -5743
rect -67 -5847 -34 -5814
rect -67 -5918 -34 -5885
rect -67 -5989 -34 -5956
rect -67 -6060 -34 -6027
rect -67 -6131 -34 -6098
rect -67 -6202 -34 -6169
rect -67 -6273 -34 -6240
rect -67 -6344 -34 -6311
rect -67 -6415 -34 -6382
rect -67 -6486 -34 -6453
rect -67 -6557 -34 -6524
rect -67 -6628 -34 -6595
rect -67 -6699 -34 -6666
rect -67 -6770 -34 -6737
rect -67 -6841 -34 -6808
rect -67 -6912 -34 -6879
rect -67 -6983 -34 -6950
rect -67 -7054 -34 -7021
rect -67 -7125 -34 -7092
rect -67 -7196 -34 -7163
rect -67 -7267 -34 -7234
rect -67 -7338 -34 -7305
rect -67 -7409 -34 -7376
rect -67 -7480 -34 -7447
rect -67 -7551 -34 -7518
rect -67 -7622 -34 -7589
rect -67 -7693 -34 -7660
rect -67 -7764 -34 -7731
rect -67 -7835 -34 -7802
rect -67 -7906 -34 -7873
rect -67 -7977 -34 -7944
rect -67 -8048 -34 -8015
rect -67 -8119 -34 -8086
rect -67 -8190 -34 -8157
rect -67 -8261 -34 -8228
rect -67 -8332 -34 -8299
rect -67 -8403 -34 -8370
rect -67 -8474 -34 -8441
rect -67 -8545 -34 -8512
rect -67 -8616 -34 -8583
rect -67 -8687 -34 -8654
rect -67 -8758 -34 -8725
rect -67 -8829 -34 -8796
rect -67 -8900 -34 -8867
rect -67 -8971 -34 -8938
rect -67 -9042 -34 -9009
rect -67 -9113 -34 -9080
rect -67 -9184 -34 -9151
rect -67 -9255 -34 -9222
rect -67 -9326 -34 -9293
rect -67 -9397 -34 -9364
rect -67 -9468 -34 -9435
rect -67 -9539 -34 -9506
rect -67 -9610 -34 -9577
rect -67 -9681 -34 -9648
rect -67 -9752 -34 -9719
rect -67 -9823 -34 -9790
rect -67 -9894 -34 -9861
rect -67 -9965 -34 -9932
rect -67 -10036 -34 -10003
rect -67 -10107 -34 -10074
rect -67 -10178 -34 -10145
rect -67 -10249 -34 -10216
rect -67 -10320 -34 -10287
rect -67 -10391 -34 -10358
rect -67 -10462 -34 -10429
rect -67 -10533 -34 -10500
rect -67 -10604 -34 -10571
rect -67 -10675 -34 -10642
rect -67 -10746 -34 -10713
rect -67 -10817 -34 -10784
rect -67 -10888 -34 -10855
rect -67 -10959 -34 -10926
rect -67 -11030 -34 -10997
rect -67 -11101 -34 -11068
rect -67 -11172 -34 -11139
rect -67 -11243 -34 -11210
rect -67 -11314 -34 -11281
rect -67 -11385 -34 -11352
rect -67 -11456 -34 -11423
rect -67 -11527 -34 -11494
rect -67 -11598 -34 -11565
rect -67 -11669 -34 -11636
rect -67 -11740 -34 -11707
rect -67 -11811 -34 -11778
rect -67 -11882 -34 -11849
rect -67 -11953 -34 -11920
rect -67 -12024 -34 -11991
rect -67 -12095 -34 -12062
rect -67 -12166 -34 -12133
rect -67 -12237 -34 -12204
rect -67 -12308 -34 -12275
rect -67 -12379 -34 -12346
rect -67 -12450 -34 -12417
rect -67 -12521 -34 -12488
rect -67 -12592 -34 -12559
rect -67 -12663 -34 -12630
rect -67 -12734 -34 -12701
rect -67 -12805 -34 -12772
rect -67 -12876 -34 -12843
rect -67 -12947 -34 -12914
rect -67 -13018 -34 -12985
rect -67 -13089 -34 -13056
rect -67 -13160 -34 -13127
rect -67 -13231 -34 -13198
rect -67 -13302 -34 -13269
rect -67 -13373 -34 -13340
rect -67 -13444 -34 -13411
rect -67 -13515 -34 -13482
rect -67 -13586 -34 -13553
rect -67 -13657 -34 -13624
rect -67 -13728 -34 -13695
rect -67 -13799 -34 -13766
rect -67 -13870 -34 -13837
rect -67 -13941 -34 -13908
rect -67 -14012 -34 -13979
rect -67 -14083 -34 -14050
rect -67 -14154 -34 -14121
rect -67 -14225 -34 -14192
rect -67 -14296 -34 -14263
rect -67 -14367 -34 -14334
rect -67 -14438 -34 -14405
rect -67 -14509 -34 -14476
rect -67 -14580 -34 -14547
rect -67 -14651 -34 -14618
rect -67 -14722 -34 -14689
rect -67 -14793 -34 -14760
rect -67 -14864 -34 -14831
rect -67 -14935 -34 -14902
rect -67 -15006 -34 -14973
rect -67 -15077 -34 -15044
rect -67 -15148 -34 -15115
rect -67 -15219 -34 -15186
rect -67 -15290 -34 -15257
rect -67 -15361 -34 -15328
rect -67 -15432 -34 -15399
rect -67 -15503 -34 -15470
rect -67 -15574 -34 -15541
rect -67 -15645 -34 -15612
rect -67 -15716 -34 -15683
rect -67 -15787 -34 -15754
rect -67 -15858 -34 -15825
rect -67 -15929 -34 -15896
rect -67 -16000 -34 -15967
rect -67 -16071 -34 -16038
rect -67 -16142 -34 -16109
rect -67 -16213 -34 -16180
rect -67 -16284 -34 -16251
rect -67 -16355 -34 -16322
rect -67 -16426 -34 -16393
rect -67 -16497 -34 -16464
rect -67 -16568 -34 -16535
rect -67 -16639 -34 -16606
rect -67 -16710 -34 -16677
rect -67 -16781 -34 -16748
rect -67 -16852 -34 -16819
rect -67 -16923 -34 -16890
rect -67 -16994 -34 -16961
rect -67 -17065 -34 -17032
rect -67 -17136 -34 -17103
rect -67 -17207 -34 -17174
rect -67 -17278 -34 -17245
rect -67 -17349 -34 -17316
rect -67 -17420 -34 -17387
rect -67 -17491 -34 -17458
rect -67 -17562 -34 -17529
rect -67 -17633 -34 -17600
rect -67 -17704 -34 -17671
rect -67 -17775 -34 -17742
rect -67 -17846 -34 -17813
rect -67 -17917 -34 -17884
rect -67 -17988 -34 -17955
rect -67 -18059 -34 -18026
rect -67 -18130 -34 -18097
rect -67 -18201 -34 -18168
rect -67 -18272 -34 -18239
rect -67 -18343 -34 -18310
rect -67 -18414 -34 -18381
rect -67 -18485 -34 -18452
rect -67 -18556 -34 -18523
rect -67 -18627 -34 -18594
rect -67 -18698 -34 -18665
rect -67 -18769 -34 -18736
rect -67 -18840 -34 -18807
rect -67 -18911 -34 -18878
rect -67 -18982 -34 -18949
rect -67 -19053 -34 -19020
rect -67 -19124 -34 -19091
rect -67 -19195 -34 -19162
rect -67 -19266 -34 -19233
rect -67 -19337 -34 -19304
rect -67 -19408 -34 -19375
rect -67 -19479 -34 -19446
rect -67 -19550 -34 -19517
rect -67 -19621 -34 -19588
rect -67 -19692 -34 -19659
rect -67 -19763 -34 -19730
rect -67 -19834 -34 -19801
rect -67 -19905 -34 -19872
rect -67 -19976 -34 -19943
rect -67 -20047 -34 -20014
rect -67 -20118 -34 -20085
rect -67 -20189 -34 -20156
rect -67 -20260 -34 -20227
rect -67 -20331 -34 -20298
rect -67 -20402 -34 -20369
rect -67 -20473 -34 -20440
rect -67 -20544 -34 -20511
rect -67 -20615 -34 -20582
rect -67 -20686 -34 -20653
rect -67 -20757 -34 -20724
rect -67 -20828 -34 -20795
rect -67 -20899 -34 -20866
rect -67 -20970 -34 -20937
rect -67 -21041 -34 -21008
rect -67 -21112 -34 -21079
rect -67 -21183 -34 -21150
rect -67 -21254 -34 -21221
rect -67 -21325 -34 -21292
rect -67 -21396 -34 -21363
rect -67 -21467 -34 -21434
rect -67 -21538 -34 -21505
rect -67 -21609 -34 -21576
rect -67 -21680 -34 -21647
rect -67 -21751 -34 -21718
rect -67 -21822 -34 -21789
rect -67 -21893 -34 -21860
rect -67 -21964 -34 -21931
rect -67 -22035 -34 -22002
rect -67 -22106 -34 -22073
rect -67 -22177 -34 -22144
rect -67 -22248 -34 -22215
rect -67 -22319 -34 -22286
rect -67 -22390 -34 -22357
rect -67 -22461 -34 -22428
rect -67 -22532 -34 -22499
rect -67 -22603 -34 -22570
rect -67 -22674 -34 -22641
rect -67 -22745 -34 -22712
rect -67 -22816 -34 -22783
rect -67 -22887 -34 -22854
rect -67 -22958 -34 -22925
rect -67 -23029 -34 -22996
rect -67 -23100 -34 -23067
rect -67 -23171 -34 -23138
rect -67 -23242 -34 -23209
rect -67 -23313 -34 -23280
rect -67 -23384 -34 -23351
rect -67 -23455 -34 -23422
rect -67 -23526 -34 -23493
rect -67 -23597 -34 -23564
rect -67 -23668 -34 -23635
rect -67 -23739 -34 -23706
rect -67 -23810 -34 -23777
rect -67 -23881 -34 -23848
rect -67 -23952 -34 -23919
rect -67 -24023 -34 -23990
rect -67 -24094 -34 -24061
rect -67 -24165 -34 -24132
rect -67 -24236 -34 -24203
rect -67 -24307 -34 -24274
rect -67 -24378 -34 -24345
rect -67 -24449 -34 -24416
rect -67 -24520 -34 -24487
rect -67 -24591 -34 -24558
rect -67 -24662 -34 -24629
rect -67 -24733 -34 -24700
rect -67 -24804 -34 -24771
rect -67 -24875 -34 -24842
rect -67 -24946 -34 -24913
rect -67 -25017 -34 -24984
rect -67 -25088 -34 -25055
rect -67 -25159 -34 -25126
rect -67 -25230 -34 -25197
rect -67 -25301 -34 -25268
rect -67 -25372 -34 -25339
rect -67 -25443 -34 -25410
rect -67 -25514 -34 -25481
rect -67 -25585 -34 -25552
rect -67 -25656 -34 -25623
rect -67 -25727 -34 -25694
rect -67 -25798 -34 -25765
rect -67 -25869 -34 -25836
rect -67 -25940 -34 -25907
rect -67 -26011 -34 -25978
rect -67 -26082 -34 -26049
rect -67 -26153 -34 -26120
rect -67 -26224 -34 -26191
rect -67 -26295 -34 -26262
rect -67 -26366 -34 -26333
rect -67 -26437 -34 -26404
rect -67 -26508 -34 -26475
rect -67 -26579 -34 -26546
rect -67 -26650 -34 -26617
rect -67 -26721 -34 -26688
rect -67 -26792 -34 -26759
rect -67 -26863 -34 -26830
rect -67 -26934 -34 -26901
rect -67 -27005 -34 -26972
rect -67 -27076 -34 -27043
rect -67 -27147 -34 -27114
rect -67 -27218 -34 -27185
rect -67 -27289 -34 -27256
rect -67 -27360 -34 -27327
rect -67 -27431 -34 -27398
rect -67 -27502 -34 -27469
rect -67 -27573 -34 -27540
rect -67 -27644 -34 -27611
rect -67 -27715 -34 -27682
rect -67 -27786 -34 -27753
rect -67 -27857 -34 -27824
rect -67 -27928 -34 -27895
rect -67 -27999 -34 -27966
rect -67 -28070 -34 -28037
rect -67 -28141 -34 -28108
rect -67 -28212 -34 -28179
rect -67 -28283 -34 -28250
rect -67 -28354 -34 -28321
rect -67 -28425 -34 -28392
rect -67 -28496 -34 -28463
rect -67 -28567 -34 -28534
rect -67 -28638 -34 -28605
rect -67 -28709 -34 -28676
rect -67 -28780 -34 -28747
rect -67 -28851 -34 -28818
rect -67 -28922 -34 -28889
rect -67 -28993 -34 -28960
rect -67 -29064 -34 -29031
rect -67 -29135 -34 -29102
rect -67 -29206 -34 -29173
rect -67 -29277 -34 -29244
rect -67 -29348 -34 -29315
rect -67 -29419 -34 -29386
rect -67 -29490 -34 -29457
rect -67 -29561 -34 -29528
rect -67 -29632 -34 -29599
rect -67 -29703 -34 -29670
rect -67 -29774 -34 -29741
rect -67 -29845 -34 -29812
rect -67 -29916 -34 -29883
rect -67 -29987 -34 -29954
rect -67 -30058 -34 -30025
rect -67 -30129 -34 -30096
rect -67 -30200 -34 -30167
rect -67 -30271 -34 -30238
rect -67 -30342 -34 -30309
rect -67 -30413 -34 -30380
rect -67 -30484 -34 -30451
rect -67 -30555 -34 -30522
rect -67 -30626 -34 -30593
rect -67 -30697 -34 -30664
rect -67 -30768 -34 -30735
rect -67 -30839 -34 -30806
rect -67 -30910 -34 -30877
rect -67 -30981 -34 -30948
rect -67 -31052 -34 -31019
rect -67 -31123 -34 -31090
rect -67 -31194 -34 -31161
rect -67 -31265 -34 -31232
rect -67 -31336 -34 -31303
rect -67 -31407 -34 -31374
rect -67 -31478 -34 -31445
rect -67 -31549 -34 -31516
rect -67 -31620 -34 -31587
rect -67 -31691 -34 -31658
rect -67 -31762 -34 -31729
rect -67 -31833 -34 -31800
rect -67 -31904 -34 -31871
rect -67 -31975 -34 -31942
rect -67 -32046 -34 -32013
rect -67 -32117 -34 -32084
rect -67 -32188 -34 -32155
rect -67 -32259 -34 -32226
rect -67 -32330 -34 -32297
rect -67 -32401 -34 -32368
rect -67 -32472 -34 -32439
rect -67 -32543 -34 -32510
rect -67 -32614 -34 -32581
rect -67 -32685 -34 -32652
rect -67 -32756 -34 -32723
rect -67 -32827 -34 -32794
rect -67 -32898 -34 -32865
rect -67 -32969 -34 -32936
rect -67 -33040 -34 -33007
rect -67 -33111 -34 -33078
rect -67 -33182 -34 -33149
rect -67 -33253 -34 -33220
rect -67 -33324 -34 -33291
rect -67 -33395 -34 -33362
rect -67 -33466 -34 -33433
rect -67 -33537 -34 -33504
rect -67 -33608 -34 -33575
rect -67 -33679 -34 -33646
rect -67 -33750 -34 -33717
rect -67 -33821 -34 -33788
rect -67 -33892 -34 -33859
rect -67 -33963 -34 -33930
rect -67 -34034 -34 -34001
rect -67 -34105 -34 -34072
rect -67 -34176 -34 -34143
rect -67 -34247 -34 -34214
rect -67 -34318 -34 -34285
rect -67 -34389 -34 -34356
rect -67 -34460 -34 -34427
rect -67 -34531 -34 -34498
rect -67 -34602 -34 -34569
rect -67 -34673 -34 -34640
rect -67 -34744 -34 -34711
rect -67 -34815 -34 -34782
rect -67 -34886 -34 -34853
rect -67 -34957 -34 -34924
rect -67 -35028 -34 -34995
rect -67 -35099 -34 -35066
rect -67 -35170 -34 -35137
rect -67 -35241 -34 -35208
rect -67 -35312 -34 -35279
rect -67 -35383 -34 -35350
rect -67 -35454 -34 -35421
rect -67 -35525 -34 -35492
rect -67 -35596 -34 -35563
rect -67 -35667 -34 -35634
rect -67 -35738 -34 -35705
rect -67 -35809 -34 -35776
rect -67 -35880 -34 -35847
rect -67 -35951 -34 -35918
rect -67 -36022 -34 -35989
rect -67 -36093 -34 -36060
rect -67 -36164 -34 -36131
rect -67 -36235 -34 -36202
rect -67 -36306 -34 -36273
rect -67 -36377 -34 -36344
rect -67 -36448 -34 -36415
rect -67 -36519 -34 -36486
rect -67 -36590 -34 -36557
rect -67 -36661 -34 -36628
rect -67 -36732 -34 -36699
rect -67 -36803 -34 -36770
rect -67 -36874 -34 -36841
rect -67 -36945 -34 -36912
rect -67 -37016 -34 -36983
rect -67 -37087 -34 -37054
rect -67 -37158 -34 -37125
rect -67 -37229 -34 -37196
rect -67 -37300 -34 -37267
rect -67 -37371 -34 -37338
rect -67 -37442 -34 -37409
rect -67 -37513 -34 -37480
rect -67 -37584 -34 -37551
rect -67 -37655 -34 -37622
rect -67 -37726 -34 -37693
rect -67 -37797 -34 -37764
rect -67 -37868 -34 -37835
rect -67 -37939 -34 -37906
rect -67 -38010 -34 -37977
rect -67 -38081 -34 -38048
rect -67 -38152 -34 -38119
rect -67 -38223 -34 -38190
rect -67 -38294 -34 -38261
rect -67 -38365 -34 -38332
rect -67 -38436 -34 -38403
rect -67 -38507 -34 -38474
rect -67 -38578 -34 -38545
rect -67 -38649 -34 -38616
rect -67 -38720 -34 -38687
rect -67 -38791 -34 -38758
rect -67 -38862 -34 -38829
rect -67 -38933 -34 -38900
rect -67 -39004 -34 -38971
rect -67 -39075 -34 -39042
rect -67 -39146 -34 -39113
rect -67 -39217 -34 -39184
rect -67 -39288 -34 -39255
rect -67 -39359 -34 -39326
rect -67 -39430 -34 -39397
rect -67 -39501 -34 -39468
rect -67 -39572 -34 -39539
rect -67 -39643 -34 -39610
rect -67 -39714 -34 -39681
rect -67 -39785 -34 -39752
rect -67 -39856 -34 -39823
rect -67 -39927 -34 -39894
rect -67 -39998 -34 -39965
rect -67 -40069 -34 -40036
rect -67 -40140 -34 -40107
rect -67 -40211 -34 -40178
rect -67 -40282 -34 -40249
rect -67 -40353 -34 -40320
rect -67 -40424 -34 -40391
rect -67 -40495 -34 -40462
rect -67 -40566 -34 -40533
rect -67 -40637 -34 -40604
rect -67 -40708 -34 -40675
rect -67 -40779 -34 -40746
rect -67 -40850 -34 -40817
rect -67 -40921 -34 -40888
rect -67 -40992 -34 -40959
rect -67 -41063 -34 -41030
rect -67 -41134 -34 -41101
rect -67 -41205 -34 -41172
rect -67 -41276 -34 -41243
rect -67 -41347 -34 -41314
rect -67 -41418 -34 -41385
rect -67 -41489 -34 -41456
rect -67 -41560 -34 -41527
rect -67 -41631 -34 -41598
rect -67 -41702 -34 -41669
rect -67 -41773 -34 -41740
rect -67 -41844 -34 -41811
rect -67 -41915 -34 -41882
rect -67 -41986 -34 -41953
rect -67 -42057 -34 -42024
rect -67 -42128 -34 -42095
rect -67 -42199 -34 -42166
rect -67 -42270 -34 -42237
rect -67 -42341 -34 -42308
rect -67 -42412 -34 -42379
rect -67 -42483 -34 -42450
rect -67 -42554 -34 -42521
rect -67 -42625 -34 -42592
rect -67 -42696 -34 -42663
rect -67 -42767 -34 -42734
rect -67 -42838 -34 -42805
rect -67 -42909 -34 -42876
rect -67 -42980 -34 -42947
rect -67 -43051 -34 -43018
rect -67 -43122 -34 -43089
rect -67 -43193 -34 -43160
rect -67 -43264 -34 -43231
rect -67 -43335 -34 -43302
rect -67 -43406 -34 -43373
rect -67 -43477 -34 -43444
rect -67 -43548 -34 -43515
rect -67 -43619 -34 -43586
rect -67 -43690 -34 -43657
rect -67 -43761 -34 -43728
rect -67 -43832 -34 -43799
rect -67 -43903 -34 -43870
rect -67 -43974 -34 -43941
rect -67 -44045 -34 -44012
rect -67 -44116 -34 -44083
rect -67 -44187 -34 -44154
rect -67 -44258 -34 -44225
rect -67 -44329 -34 -44296
rect -67 -44400 -34 -44367
rect -67 -44471 -34 -44438
rect -67 -44542 -34 -44509
rect -67 -44613 -34 -44580
rect -67 -44684 -34 -44651
rect -67 -44755 -34 -44722
rect -67 -44826 -34 -44793
rect -67 -44897 -34 -44864
rect -67 -44968 -34 -44935
rect -67 -45039 -34 -45006
rect -67 -45110 -34 -45077
rect -67 -45181 -34 -45148
rect -67 -45252 -34 -45219
rect -67 -45323 -34 -45290
rect -67 -45394 -34 -45361
rect -67 -45465 -34 -45432
rect -67 -45536 -34 -45503
rect -67 -45607 -34 -45574
rect -67 -45678 -34 -45645
rect -67 -45749 -34 -45716
rect -67 -45820 -34 -45787
rect -67 -45891 -34 -45858
rect -67 -45962 -34 -45929
rect -67 -46033 -34 -46000
rect -67 -46104 -34 -46071
rect -67 -46175 -34 -46142
rect -67 -46246 -34 -46213
rect -67 -46317 -34 -46284
rect -67 -46388 -34 -46355
rect -67 -46459 -34 -46426
rect -67 -46530 -34 -46497
rect -67 -46601 -34 -46568
rect -67 -46672 -34 -46639
rect -67 -46743 -34 -46710
rect -67 -46814 -34 -46781
rect -67 -46885 -34 -46852
rect -67 -46956 -34 -46923
rect -67 -47027 -34 -46994
rect -67 -47098 -34 -47065
rect -67 -47169 -34 -47136
rect -67 -47240 -34 -47207
rect -67 -47311 -34 -47278
rect -67 -47382 -34 -47349
rect -67 -47453 -34 -47420
rect -67 -47524 -34 -47491
rect -67 -47595 -34 -47562
rect -67 -47666 -34 -47633
rect -67 -47737 -34 -47704
rect -67 -47808 -34 -47775
rect -67 -47879 -34 -47846
rect -67 -47950 -34 -47917
rect -67 -48021 -34 -47988
rect -67 -48092 -34 -48059
rect -67 -48163 -34 -48130
rect -67 -48234 -34 -48201
rect -67 -48305 -34 -48272
rect -67 -48376 -34 -48343
rect -67 -48447 -34 -48414
rect -67 -48518 -34 -48485
rect -67 -48589 -34 -48556
rect -67 -48660 -34 -48627
rect -67 -48731 -34 -48698
rect -67 -48802 -34 -48769
rect -67 -48873 -34 -48840
rect -67 -48944 -34 -48911
rect -67 -49015 -34 -48982
rect -67 -49086 -34 -49053
rect -67 -49157 -34 -49124
rect -67 -49228 -34 -49195
rect -67 -49299 -34 -49266
rect -67 -49370 -34 -49337
rect -67 -49441 -34 -49408
rect -67 -49512 -34 -49479
rect -67 -49583 -34 -49550
rect -67 -49654 -34 -49621
rect -67 -49725 -34 -49692
rect -67 -49796 -34 -49763
rect -67 -49867 -34 -49834
rect -67 -49938 -34 -49905
rect -67 -50009 -34 -49976
rect -67 -50080 -34 -50047
rect -67 -50151 -34 -50118
rect -67 -50222 -34 -50189
rect -67 -50293 -34 -50260
rect -67 -50364 -34 -50331
rect -67 -50435 -34 -50402
rect -67 -50506 -34 -50473
rect -67 -50577 -34 -50544
rect -67 -50648 -34 -50615
rect -67 -50719 -34 -50686
rect -67 -50790 -34 -50757
rect -67 -50861 -34 -50828
rect -67 -50932 -34 -50899
rect -67 -51003 -34 -50970
rect -67 -51074 -34 -51041
rect -67 -51145 -34 -51112
rect -67 -51216 -34 -51183
rect -67 -51287 -34 -51254
rect -67 -51358 -34 -51325
rect -67 -51429 -34 -51396
rect -67 -51500 -34 -51467
rect -67 -51571 -34 -51538
rect -67 -51642 -34 -51609
rect -67 -51713 -34 -51680
rect -67 -51784 -34 -51751
rect -67 -51855 -34 -51822
rect -67 -51926 -34 -51893
rect -67 -51997 -34 -51964
rect -67 -52068 -34 -52035
rect -67 -52139 -34 -52106
rect -67 -52210 -34 -52177
rect -67 -52281 -34 -52248
rect -67 -52352 -34 -52319
rect -67 -52423 -34 -52390
rect -67 -52494 -34 -52461
rect -67 -52565 -34 -52532
rect -67 -52636 -34 -52603
rect -67 -52707 -34 -52674
rect -67 -52778 -34 -52745
rect -67 -52849 -34 -52816
rect -67 -52920 -34 -52887
rect -67 -52991 -34 -52958
rect -67 -53062 -34 -53029
rect -67 -53133 -34 -53100
rect -67 -53204 -34 -53171
rect -67 -53275 -34 -53242
rect -67 -53346 -34 -53313
rect -67 -53417 -34 -53384
rect -67 -53488 -34 -53455
rect -67 -53559 -34 -53526
rect -67 -53630 -34 -53597
rect -67 -53701 -34 -53668
rect -67 -53772 -34 -53739
rect -67 -53843 -34 -53810
rect -67 -53914 -34 -53881
rect -67 -53985 -34 -53952
rect -67 -54056 -34 -54023
rect -67 -54127 -34 -54094
rect -67 -54198 -34 -54165
rect -67 -54269 -34 -54236
rect -67 -54340 -34 -54307
rect -67 -54411 -34 -54378
rect -67 -54482 -34 -54449
rect -67 -54553 -34 -54520
rect -67 -54624 -34 -54591
rect -67 -54695 -34 -54662
rect -67 -54766 -34 -54733
rect -67 -54837 -34 -54804
rect -67 -54908 -34 -54875
rect -67 -54979 -34 -54946
rect -67 -55050 -34 -55017
rect -67 -55121 -34 -55088
rect -67 -55192 -34 -55159
rect -67 -55263 -34 -55230
rect -67 -55334 -34 -55301
rect -67 -55405 -34 -55372
rect -67 -55476 -34 -55443
rect -67 -55547 -34 -55514
rect -67 -55618 -34 -55585
rect -67 -55689 -34 -55656
rect -67 -55760 -34 -55727
rect -67 -55831 -34 -55798
rect -67 -55902 -34 -55869
rect -67 -55973 -34 -55940
rect -67 -56044 -34 -56011
rect -67 -56115 -34 -56082
rect -67 -56186 -34 -56153
rect -67 -56257 -34 -56224
rect -67 -56328 -34 -56295
rect -67 -56399 -34 -56366
rect -67 -56470 -34 -56437
rect -67 -56541 -34 -56508
rect -67 -56612 -34 -56579
rect -67 -56683 -34 -56650
rect -67 -56754 -34 -56721
rect -67 -56825 -34 -56792
rect -67 -56896 -34 -56863
rect -67 -56967 -34 -56934
rect -67 -57038 -34 -57005
rect -67 -57109 -34 -57076
rect -67 -57180 -34 -57147
rect -67 -57251 -34 -57218
rect -67 -57322 -34 -57289
rect -67 -57393 -34 -57360
rect -67 -57464 -34 -57431
rect -67 -57535 -34 -57502
rect -67 -57606 -34 -57573
rect -67 -57677 -34 -57644
rect -67 -57748 -34 -57715
rect -67 -57819 -34 -57786
rect -67 -57890 -34 -57857
rect -67 -57961 -34 -57928
rect -67 -58032 -34 -57999
rect -67 -58103 -34 -58070
rect -67 -58174 -34 -58141
rect -67 -58245 -34 -58212
rect -67 -58316 -34 -58283
rect -67 -58387 -34 -58354
rect -67 -58458 -34 -58425
rect -67 -58529 -34 -58496
rect -67 -58600 -34 -58567
rect -67 -58671 -34 -58638
rect -67 -58742 -34 -58709
rect -67 -58813 -34 -58780
rect -67 -58884 -34 -58851
rect -67 -58955 -34 -58922
rect -67 -59026 -34 -58993
rect -67 -59097 -34 -59064
rect -67 -59168 -34 -59135
rect -67 -59239 -34 -59206
rect -67 -59310 -34 -59277
rect -67 -59381 -34 -59348
rect -67 -59452 -34 -59419
rect -67 -59523 -34 -59490
rect -67 -59594 -34 -59561
rect -67 -59665 -34 -59632
rect -67 -59736 -34 -59703
rect -67 -59807 -34 -59774
rect -67 -59878 -34 -59845
rect -67 -59949 -34 -59916
rect -67 -60020 -34 -59987
rect -67 -60091 -34 -60058
rect -67 -60162 -34 -60129
rect -67 -60233 -34 -60200
rect -67 -60304 -34 -60271
rect -67 -60375 -34 -60342
rect -67 -60446 -34 -60413
rect -67 -60517 -34 -60484
rect -67 -60588 -34 -60555
rect -67 -60659 -34 -60626
rect -67 -60730 -34 -60697
rect -67 -60801 -34 -60768
rect -67 -60872 -34 -60839
rect -67 -60943 -34 -60910
rect -67 -61014 -34 -60981
rect -67 -61085 -34 -61052
rect -67 -61156 -34 -61123
rect -67 -61227 -34 -61194
rect -67 -61298 -34 -61265
rect -67 -61369 -34 -61336
rect -67 -61440 -34 -61407
rect -67 -61511 -34 -61478
rect -67 -61582 -34 -61549
rect -67 -61653 -34 -61620
rect -67 -61724 -34 -61691
rect -67 -61795 -34 -61762
rect -67 -61866 -34 -61833
rect -67 -61937 -34 -61904
rect -67 -62008 -34 -61975
rect -67 -62079 -34 -62046
rect -67 -62150 -34 -62117
rect -67 -62221 -34 -62188
rect -67 -62292 -34 -62259
rect -67 -62363 -34 -62330
rect -67 -62434 -34 -62401
rect -67 -62505 -34 -62472
rect -67 -62576 -34 -62543
rect -67 -62647 -34 -62614
rect -67 -62718 -34 -62685
rect -67 -62789 -34 -62756
rect -67 -62860 -34 -62827
rect -67 -62931 -34 -62898
rect -67 -63002 -34 -62969
rect -67 -63073 -34 -63040
rect -67 -63144 -34 -63111
rect -67 -63215 -34 -63182
rect -67 -63286 -34 -63253
rect -67 -63357 -34 -63324
rect -67 -63428 -34 -63395
rect -67 -63499 -34 -63466
rect -67 -63570 -34 -63537
rect -67 -63641 -34 -63608
rect -67 -63712 -34 -63679
rect -67 -63783 -34 -63750
rect -67 -63854 -34 -63821
rect -67 -63925 -34 -63892
rect -67 -63996 -34 -63963
rect -67 -64067 -34 -64034
rect -67 -64138 -34 -64105
rect -67 -64209 -34 -64176
rect -67 -64280 -34 -64247
rect -67 -64351 -34 -64318
rect -67 -64422 -34 -64389
rect -67 -64493 -34 -64460
rect -67 -64564 -34 -64531
rect -67 -64635 -34 -64602
rect -67 -64706 -34 -64673
rect -67 -64777 -34 -64744
rect -67 -64848 -34 -64815
rect -67 -64919 -34 -64886
rect -67 -64990 -34 -64957
rect -67 -65061 -34 -65028
rect -67 -65132 -34 -65099
rect -67 -65203 -34 -65170
rect -67 -65274 -34 -65241
rect -67 -65345 -34 -65312
rect -67 -65416 -34 -65383
rect -67 -65487 -34 -65454
rect -67 -65558 -34 -65525
rect -67 -65629 -34 -65596
rect -67 -65700 -34 -65667
rect -67 -65771 -34 -65738
rect -67 -65842 -34 -65809
rect -67 -65913 -34 -65880
rect -67 -65984 -34 -65951
rect -67 -66055 -34 -66022
rect -67 -66126 -34 -66093
rect -67 -66197 -34 -66164
rect -67 -66268 -34 -66235
rect -67 -66339 -34 -66306
rect -67 -66410 -34 -66377
rect -67 -66481 -34 -66448
rect -67 -66552 -34 -66519
rect -67 -66623 -34 -66590
rect -67 -66694 -34 -66661
rect -67 -66765 -34 -66732
rect -67 -66836 -34 -66803
rect -67 -66907 -34 -66874
rect -67 -66978 -34 -66945
rect -67 -67049 -34 -67016
rect -67 -67120 -34 -67087
rect -67 -67191 -34 -67158
rect -67 -67262 -34 -67229
rect -67 -67333 -34 -67300
rect -67 -67404 -34 -67371
rect -67 -67475 -34 -67442
rect -67 -67546 -34 -67513
rect -67 -67617 -34 -67584
rect -67 -67688 -34 -67655
rect -67 -67759 -34 -67726
rect -67 -67830 -34 -67797
rect -67 -67901 -34 -67868
rect -67 -67972 -34 -67939
rect -67 -68043 -34 -68010
rect -67 -68114 -34 -68081
rect -67 -68185 -34 -68152
rect -67 -68256 -34 -68223
rect -67 -68327 -34 -68294
rect -67 -68398 -34 -68365
rect -67 -68469 -34 -68436
rect -67 -68540 -34 -68507
rect -67 -68611 -34 -68578
rect -67 -68682 -34 -68649
rect -67 -68753 -34 -68720
rect -67 -68824 -34 -68791
rect -67 -68895 -34 -68862
rect -67 -68966 -34 -68933
rect -67 -69037 -34 -69004
rect -67 -69108 -34 -69075
rect -67 -69179 -34 -69146
rect -67 -69250 -34 -69217
rect -67 -69321 -34 -69288
rect -67 -69392 -34 -69359
rect -67 -69463 -34 -69430
rect -67 -69534 -34 -69501
rect -67 -69605 -34 -69572
rect -67 -69676 -34 -69643
rect -67 -69747 -34 -69714
rect -67 -69818 -34 -69785
rect -67 -69889 -34 -69856
rect -67 -69960 -34 -69927
rect -67 -70031 -34 -69998
rect -67 -70102 -34 -70069
rect -67 -70173 -34 -70140
rect -67 -70244 -34 -70211
rect -67 -70315 -34 -70282
rect -67 -70386 -34 -70353
rect -67 -70457 -34 -70424
rect -67 -70528 -34 -70495
rect -67 -70599 -34 -70566
rect -67 -70670 -34 -70637
rect -67 -70741 -34 -70708
rect -67 -70812 -34 -70779
rect -67 -70883 -34 -70850
rect -67 -70954 -34 -70921
rect -67 -71025 -34 -70992
rect -67 -71096 -34 -71063
rect -67 -71167 -34 -71134
rect -67 -71238 -34 -71205
rect -67 -71309 -34 -71276
rect -67 -71380 -34 -71347
rect -67 -71451 -34 -71418
rect -67 -71522 -34 -71489
rect -67 -71593 -34 -71560
rect -67 -71664 -34 -71631
rect -67 -71735 -34 -71702
rect -67 -71806 -34 -71773
rect -67 -71877 -34 -71844
rect -67 -71948 -34 -71915
rect -67 -72019 -34 -71986
rect -67 -72090 -34 -72057
rect -67 -72161 -34 -72128
rect -67 -72232 -34 -72199
rect -67 -72303 -34 -72270
rect -67 -72374 -34 -72341
rect -67 -72445 -34 -72412
rect -67 -72516 -34 -72483
rect -67 -72587 -34 -72554
rect -67 -72658 -34 -72625
rect 0 -72704 33 41
rect 0 -72737 33 -72704
rect 83 -72704 116 41
rect 166 -72704 199 41
rect 166 -72737 199 -72704
rect 249 -72704 282 41
rect 249 -72737 282 -72704
rect 332 -72704 365 41
rect 415 -72704 448 41
rect 415 -72737 448 -72704
rect 498 -72704 531 41
rect 498 -72737 531 -72704
rect 581 -72704 614 41
rect 664 -72704 697 41
rect 664 -72737 697 -72704
rect 747 -72704 780 41
rect 747 -72737 780 -72704
rect 830 -72704 863 41
rect 913 -72704 946 41
rect 913 -72737 946 -72704
rect 913 19 946 52
rect 913 138 946 171
rect 904 194 955 227
rect 904 227 955 244
rect 747 19 780 52
rect 747 138 780 171
rect 738 194 789 227
rect 738 227 789 244
rect 664 19 697 52
rect 664 138 697 171
rect 655 194 706 227
rect 655 227 706 244
rect 498 19 531 52
rect 498 138 531 171
rect 489 194 540 227
rect 489 227 540 244
rect 415 19 448 52
rect 415 138 448 171
rect 406 194 457 227
rect 406 227 457 244
rect 249 19 282 52
rect 249 138 282 171
rect 240 194 291 227
rect 240 227 291 244
rect 166 19 199 52
rect 166 138 199 171
rect 157 194 208 227
rect 157 227 208 244
rect 0 19 33 52
rect 0 138 33 171
rect -9 194 42 227
rect -9 227 42 244
rect -27 69 973 117
rect -60 69 -27 199
rect 830 41 863 69
rect 581 41 614 69
rect 332 41 365 69
rect 83 41 116 69
rect -25 244 971 292
<< viali >>
rect 921 27 938 44
rect 921 146 938 163
rect 755 27 772 44
rect 755 146 772 163
rect 672 27 689 44
rect 672 146 689 163
rect 506 27 523 44
rect 506 146 523 163
rect 423 27 440 44
rect 423 146 440 163
rect 257 27 274 44
rect 257 146 274 163
rect 174 27 191 44
rect 174 146 191 163
rect 8 27 25 44
rect 8 146 25 163
<< metal1 >>
rect 913 19 946 171
rect 747 19 780 171
rect 664 19 697 171
rect 498 19 531 171
rect 415 19 448 171
rect 249 19 282 171
rect 166 19 199 171
rect 0 19 33 171
<< labels >>
flabel locali -67 -25 -34 8 0 FreeSerif 160 0 0 0 word0
port 100 nsew
flabel locali -67 -96 -34 -63 0 FreeSerif 160 0 0 0 word1
port 101 nsew
flabel locali -67 -167 -34 -134 0 FreeSerif 160 0 0 0 word2
port 102 nsew
flabel locali -67 -238 -34 -205 0 FreeSerif 160 0 0 0 word3
port 103 nsew
flabel locali -67 -309 -34 -276 0 FreeSerif 160 0 0 0 word4
port 104 nsew
flabel locali -67 -380 -34 -347 0 FreeSerif 160 0 0 0 word5
port 105 nsew
flabel locali -67 -451 -34 -418 0 FreeSerif 160 0 0 0 word6
port 106 nsew
flabel locali -67 -522 -34 -489 0 FreeSerif 160 0 0 0 word7
port 107 nsew
flabel locali -67 -593 -34 -560 0 FreeSerif 160 0 0 0 word8
port 108 nsew
flabel locali -67 -664 -34 -631 0 FreeSerif 160 0 0 0 word9
port 109 nsew
flabel locali -67 -735 -34 -702 0 FreeSerif 160 0 0 0 word10
port 110 nsew
flabel locali -67 -806 -34 -773 0 FreeSerif 160 0 0 0 word11
port 111 nsew
flabel locali -67 -877 -34 -844 0 FreeSerif 160 0 0 0 word12
port 112 nsew
flabel locali -67 -948 -34 -915 0 FreeSerif 160 0 0 0 word13
port 113 nsew
flabel locali -67 -1019 -34 -986 0 FreeSerif 160 0 0 0 word14
port 114 nsew
flabel locali -67 -1090 -34 -1057 0 FreeSerif 160 0 0 0 word15
port 115 nsew
flabel locali -67 -1161 -34 -1128 0 FreeSerif 160 0 0 0 word16
port 116 nsew
flabel locali -67 -1232 -34 -1199 0 FreeSerif 160 0 0 0 word17
port 117 nsew
flabel locali -67 -1303 -34 -1270 0 FreeSerif 160 0 0 0 word18
port 118 nsew
flabel locali -67 -1374 -34 -1341 0 FreeSerif 160 0 0 0 word19
port 119 nsew
flabel locali -67 -1445 -34 -1412 0 FreeSerif 160 0 0 0 word20
port 120 nsew
flabel locali -67 -1516 -34 -1483 0 FreeSerif 160 0 0 0 word21
port 121 nsew
flabel locali -67 -1587 -34 -1554 0 FreeSerif 160 0 0 0 word22
port 122 nsew
flabel locali -67 -1658 -34 -1625 0 FreeSerif 160 0 0 0 word23
port 123 nsew
flabel locali -67 -1729 -34 -1696 0 FreeSerif 160 0 0 0 word24
port 124 nsew
flabel locali -67 -1800 -34 -1767 0 FreeSerif 160 0 0 0 word25
port 125 nsew
flabel locali -67 -1871 -34 -1838 0 FreeSerif 160 0 0 0 word26
port 126 nsew
flabel locali -67 -1942 -34 -1909 0 FreeSerif 160 0 0 0 word27
port 127 nsew
flabel locali -67 -2013 -34 -1980 0 FreeSerif 160 0 0 0 word28
port 128 nsew
flabel locali -67 -2084 -34 -2051 0 FreeSerif 160 0 0 0 word29
port 129 nsew
flabel locali -67 -2155 -34 -2122 0 FreeSerif 160 0 0 0 word30
port 130 nsew
flabel locali -67 -2226 -34 -2193 0 FreeSerif 160 0 0 0 word31
port 131 nsew
flabel locali -67 -2297 -34 -2264 0 FreeSerif 160 0 0 0 word32
port 132 nsew
flabel locali -67 -2368 -34 -2335 0 FreeSerif 160 0 0 0 word33
port 133 nsew
flabel locali -67 -2439 -34 -2406 0 FreeSerif 160 0 0 0 word34
port 134 nsew
flabel locali -67 -2510 -34 -2477 0 FreeSerif 160 0 0 0 word35
port 135 nsew
flabel locali -67 -2581 -34 -2548 0 FreeSerif 160 0 0 0 word36
port 136 nsew
flabel locali -67 -2652 -34 -2619 0 FreeSerif 160 0 0 0 word37
port 137 nsew
flabel locali -67 -2723 -34 -2690 0 FreeSerif 160 0 0 0 word38
port 138 nsew
flabel locali -67 -2794 -34 -2761 0 FreeSerif 160 0 0 0 word39
port 139 nsew
flabel locali -67 -2865 -34 -2832 0 FreeSerif 160 0 0 0 word40
port 140 nsew
flabel locali -67 -2936 -34 -2903 0 FreeSerif 160 0 0 0 word41
port 141 nsew
flabel locali -67 -3007 -34 -2974 0 FreeSerif 160 0 0 0 word42
port 142 nsew
flabel locali -67 -3078 -34 -3045 0 FreeSerif 160 0 0 0 word43
port 143 nsew
flabel locali -67 -3149 -34 -3116 0 FreeSerif 160 0 0 0 word44
port 144 nsew
flabel locali -67 -3220 -34 -3187 0 FreeSerif 160 0 0 0 word45
port 145 nsew
flabel locali -67 -3291 -34 -3258 0 FreeSerif 160 0 0 0 word46
port 146 nsew
flabel locali -67 -3362 -34 -3329 0 FreeSerif 160 0 0 0 word47
port 147 nsew
flabel locali -67 -3433 -34 -3400 0 FreeSerif 160 0 0 0 word48
port 148 nsew
flabel locali -67 -3504 -34 -3471 0 FreeSerif 160 0 0 0 word49
port 149 nsew
flabel locali -67 -3575 -34 -3542 0 FreeSerif 160 0 0 0 word50
port 150 nsew
flabel locali -67 -3646 -34 -3613 0 FreeSerif 160 0 0 0 word51
port 151 nsew
flabel locali -67 -3717 -34 -3684 0 FreeSerif 160 0 0 0 word52
port 152 nsew
flabel locali -67 -3788 -34 -3755 0 FreeSerif 160 0 0 0 word53
port 153 nsew
flabel locali -67 -3859 -34 -3826 0 FreeSerif 160 0 0 0 word54
port 154 nsew
flabel locali -67 -3930 -34 -3897 0 FreeSerif 160 0 0 0 word55
port 155 nsew
flabel locali -67 -4001 -34 -3968 0 FreeSerif 160 0 0 0 word56
port 156 nsew
flabel locali -67 -4072 -34 -4039 0 FreeSerif 160 0 0 0 word57
port 157 nsew
flabel locali -67 -4143 -34 -4110 0 FreeSerif 160 0 0 0 word58
port 158 nsew
flabel locali -67 -4214 -34 -4181 0 FreeSerif 160 0 0 0 word59
port 159 nsew
flabel locali -67 -4285 -34 -4252 0 FreeSerif 160 0 0 0 word60
port 160 nsew
flabel locali -67 -4356 -34 -4323 0 FreeSerif 160 0 0 0 word61
port 161 nsew
flabel locali -67 -4427 -34 -4394 0 FreeSerif 160 0 0 0 word62
port 162 nsew
flabel locali -67 -4498 -34 -4465 0 FreeSerif 160 0 0 0 word63
port 163 nsew
flabel locali -67 -4569 -34 -4536 0 FreeSerif 160 0 0 0 word64
port 164 nsew
flabel locali -67 -4640 -34 -4607 0 FreeSerif 160 0 0 0 word65
port 165 nsew
flabel locali -67 -4711 -34 -4678 0 FreeSerif 160 0 0 0 word66
port 166 nsew
flabel locali -67 -4782 -34 -4749 0 FreeSerif 160 0 0 0 word67
port 167 nsew
flabel locali -67 -4853 -34 -4820 0 FreeSerif 160 0 0 0 word68
port 168 nsew
flabel locali -67 -4924 -34 -4891 0 FreeSerif 160 0 0 0 word69
port 169 nsew
flabel locali -67 -4995 -34 -4962 0 FreeSerif 160 0 0 0 word70
port 170 nsew
flabel locali -67 -5066 -34 -5033 0 FreeSerif 160 0 0 0 word71
port 171 nsew
flabel locali -67 -5137 -34 -5104 0 FreeSerif 160 0 0 0 word72
port 172 nsew
flabel locali -67 -5208 -34 -5175 0 FreeSerif 160 0 0 0 word73
port 173 nsew
flabel locali -67 -5279 -34 -5246 0 FreeSerif 160 0 0 0 word74
port 174 nsew
flabel locali -67 -5350 -34 -5317 0 FreeSerif 160 0 0 0 word75
port 175 nsew
flabel locali -67 -5421 -34 -5388 0 FreeSerif 160 0 0 0 word76
port 176 nsew
flabel locali -67 -5492 -34 -5459 0 FreeSerif 160 0 0 0 word77
port 177 nsew
flabel locali -67 -5563 -34 -5530 0 FreeSerif 160 0 0 0 word78
port 178 nsew
flabel locali -67 -5634 -34 -5601 0 FreeSerif 160 0 0 0 word79
port 179 nsew
flabel locali -67 -5705 -34 -5672 0 FreeSerif 160 0 0 0 word80
port 180 nsew
flabel locali -67 -5776 -34 -5743 0 FreeSerif 160 0 0 0 word81
port 181 nsew
flabel locali -67 -5847 -34 -5814 0 FreeSerif 160 0 0 0 word82
port 182 nsew
flabel locali -67 -5918 -34 -5885 0 FreeSerif 160 0 0 0 word83
port 183 nsew
flabel locali -67 -5989 -34 -5956 0 FreeSerif 160 0 0 0 word84
port 184 nsew
flabel locali -67 -6060 -34 -6027 0 FreeSerif 160 0 0 0 word85
port 185 nsew
flabel locali -67 -6131 -34 -6098 0 FreeSerif 160 0 0 0 word86
port 186 nsew
flabel locali -67 -6202 -34 -6169 0 FreeSerif 160 0 0 0 word87
port 187 nsew
flabel locali -67 -6273 -34 -6240 0 FreeSerif 160 0 0 0 word88
port 188 nsew
flabel locali -67 -6344 -34 -6311 0 FreeSerif 160 0 0 0 word89
port 189 nsew
flabel locali -67 -6415 -34 -6382 0 FreeSerif 160 0 0 0 word90
port 190 nsew
flabel locali -67 -6486 -34 -6453 0 FreeSerif 160 0 0 0 word91
port 191 nsew
flabel locali -67 -6557 -34 -6524 0 FreeSerif 160 0 0 0 word92
port 192 nsew
flabel locali -67 -6628 -34 -6595 0 FreeSerif 160 0 0 0 word93
port 193 nsew
flabel locali -67 -6699 -34 -6666 0 FreeSerif 160 0 0 0 word94
port 194 nsew
flabel locali -67 -6770 -34 -6737 0 FreeSerif 160 0 0 0 word95
port 195 nsew
flabel locali -67 -6841 -34 -6808 0 FreeSerif 160 0 0 0 word96
port 196 nsew
flabel locali -67 -6912 -34 -6879 0 FreeSerif 160 0 0 0 word97
port 197 nsew
flabel locali -67 -6983 -34 -6950 0 FreeSerif 160 0 0 0 word98
port 198 nsew
flabel locali -67 -7054 -34 -7021 0 FreeSerif 160 0 0 0 word99
port 199 nsew
flabel locali -67 -7125 -34 -7092 0 FreeSerif 160 0 0 0 word100
port 200 nsew
flabel locali -67 -7196 -34 -7163 0 FreeSerif 160 0 0 0 word101
port 201 nsew
flabel locali -67 -7267 -34 -7234 0 FreeSerif 160 0 0 0 word102
port 202 nsew
flabel locali -67 -7338 -34 -7305 0 FreeSerif 160 0 0 0 word103
port 203 nsew
flabel locali -67 -7409 -34 -7376 0 FreeSerif 160 0 0 0 word104
port 204 nsew
flabel locali -67 -7480 -34 -7447 0 FreeSerif 160 0 0 0 word105
port 205 nsew
flabel locali -67 -7551 -34 -7518 0 FreeSerif 160 0 0 0 word106
port 206 nsew
flabel locali -67 -7622 -34 -7589 0 FreeSerif 160 0 0 0 word107
port 207 nsew
flabel locali -67 -7693 -34 -7660 0 FreeSerif 160 0 0 0 word108
port 208 nsew
flabel locali -67 -7764 -34 -7731 0 FreeSerif 160 0 0 0 word109
port 209 nsew
flabel locali -67 -7835 -34 -7802 0 FreeSerif 160 0 0 0 word110
port 210 nsew
flabel locali -67 -7906 -34 -7873 0 FreeSerif 160 0 0 0 word111
port 211 nsew
flabel locali -67 -7977 -34 -7944 0 FreeSerif 160 0 0 0 word112
port 212 nsew
flabel locali -67 -8048 -34 -8015 0 FreeSerif 160 0 0 0 word113
port 213 nsew
flabel locali -67 -8119 -34 -8086 0 FreeSerif 160 0 0 0 word114
port 214 nsew
flabel locali -67 -8190 -34 -8157 0 FreeSerif 160 0 0 0 word115
port 215 nsew
flabel locali -67 -8261 -34 -8228 0 FreeSerif 160 0 0 0 word116
port 216 nsew
flabel locali -67 -8332 -34 -8299 0 FreeSerif 160 0 0 0 word117
port 217 nsew
flabel locali -67 -8403 -34 -8370 0 FreeSerif 160 0 0 0 word118
port 218 nsew
flabel locali -67 -8474 -34 -8441 0 FreeSerif 160 0 0 0 word119
port 219 nsew
flabel locali -67 -8545 -34 -8512 0 FreeSerif 160 0 0 0 word120
port 220 nsew
flabel locali -67 -8616 -34 -8583 0 FreeSerif 160 0 0 0 word121
port 221 nsew
flabel locali -67 -8687 -34 -8654 0 FreeSerif 160 0 0 0 word122
port 222 nsew
flabel locali -67 -8758 -34 -8725 0 FreeSerif 160 0 0 0 word123
port 223 nsew
flabel locali -67 -8829 -34 -8796 0 FreeSerif 160 0 0 0 word124
port 224 nsew
flabel locali -67 -8900 -34 -8867 0 FreeSerif 160 0 0 0 word125
port 225 nsew
flabel locali -67 -8971 -34 -8938 0 FreeSerif 160 0 0 0 word126
port 226 nsew
flabel locali -67 -9042 -34 -9009 0 FreeSerif 160 0 0 0 word127
port 227 nsew
flabel locali -67 -9113 -34 -9080 0 FreeSerif 160 0 0 0 word128
port 228 nsew
flabel locali -67 -9184 -34 -9151 0 FreeSerif 160 0 0 0 word129
port 229 nsew
flabel locali -67 -9255 -34 -9222 0 FreeSerif 160 0 0 0 word130
port 230 nsew
flabel locali -67 -9326 -34 -9293 0 FreeSerif 160 0 0 0 word131
port 231 nsew
flabel locali -67 -9397 -34 -9364 0 FreeSerif 160 0 0 0 word132
port 232 nsew
flabel locali -67 -9468 -34 -9435 0 FreeSerif 160 0 0 0 word133
port 233 nsew
flabel locali -67 -9539 -34 -9506 0 FreeSerif 160 0 0 0 word134
port 234 nsew
flabel locali -67 -9610 -34 -9577 0 FreeSerif 160 0 0 0 word135
port 235 nsew
flabel locali -67 -9681 -34 -9648 0 FreeSerif 160 0 0 0 word136
port 236 nsew
flabel locali -67 -9752 -34 -9719 0 FreeSerif 160 0 0 0 word137
port 237 nsew
flabel locali -67 -9823 -34 -9790 0 FreeSerif 160 0 0 0 word138
port 238 nsew
flabel locali -67 -9894 -34 -9861 0 FreeSerif 160 0 0 0 word139
port 239 nsew
flabel locali -67 -9965 -34 -9932 0 FreeSerif 160 0 0 0 word140
port 240 nsew
flabel locali -67 -10036 -34 -10003 0 FreeSerif 160 0 0 0 word141
port 241 nsew
flabel locali -67 -10107 -34 -10074 0 FreeSerif 160 0 0 0 word142
port 242 nsew
flabel locali -67 -10178 -34 -10145 0 FreeSerif 160 0 0 0 word143
port 243 nsew
flabel locali -67 -10249 -34 -10216 0 FreeSerif 160 0 0 0 word144
port 244 nsew
flabel locali -67 -10320 -34 -10287 0 FreeSerif 160 0 0 0 word145
port 245 nsew
flabel locali -67 -10391 -34 -10358 0 FreeSerif 160 0 0 0 word146
port 246 nsew
flabel locali -67 -10462 -34 -10429 0 FreeSerif 160 0 0 0 word147
port 247 nsew
flabel locali -67 -10533 -34 -10500 0 FreeSerif 160 0 0 0 word148
port 248 nsew
flabel locali -67 -10604 -34 -10571 0 FreeSerif 160 0 0 0 word149
port 249 nsew
flabel locali -67 -10675 -34 -10642 0 FreeSerif 160 0 0 0 word150
port 250 nsew
flabel locali -67 -10746 -34 -10713 0 FreeSerif 160 0 0 0 word151
port 251 nsew
flabel locali -67 -10817 -34 -10784 0 FreeSerif 160 0 0 0 word152
port 252 nsew
flabel locali -67 -10888 -34 -10855 0 FreeSerif 160 0 0 0 word153
port 253 nsew
flabel locali -67 -10959 -34 -10926 0 FreeSerif 160 0 0 0 word154
port 254 nsew
flabel locali -67 -11030 -34 -10997 0 FreeSerif 160 0 0 0 word155
port 255 nsew
flabel locali -67 -11101 -34 -11068 0 FreeSerif 160 0 0 0 word156
port 256 nsew
flabel locali -67 -11172 -34 -11139 0 FreeSerif 160 0 0 0 word157
port 257 nsew
flabel locali -67 -11243 -34 -11210 0 FreeSerif 160 0 0 0 word158
port 258 nsew
flabel locali -67 -11314 -34 -11281 0 FreeSerif 160 0 0 0 word159
port 259 nsew
flabel locali -67 -11385 -34 -11352 0 FreeSerif 160 0 0 0 word160
port 260 nsew
flabel locali -67 -11456 -34 -11423 0 FreeSerif 160 0 0 0 word161
port 261 nsew
flabel locali -67 -11527 -34 -11494 0 FreeSerif 160 0 0 0 word162
port 262 nsew
flabel locali -67 -11598 -34 -11565 0 FreeSerif 160 0 0 0 word163
port 263 nsew
flabel locali -67 -11669 -34 -11636 0 FreeSerif 160 0 0 0 word164
port 264 nsew
flabel locali -67 -11740 -34 -11707 0 FreeSerif 160 0 0 0 word165
port 265 nsew
flabel locali -67 -11811 -34 -11778 0 FreeSerif 160 0 0 0 word166
port 266 nsew
flabel locali -67 -11882 -34 -11849 0 FreeSerif 160 0 0 0 word167
port 267 nsew
flabel locali -67 -11953 -34 -11920 0 FreeSerif 160 0 0 0 word168
port 268 nsew
flabel locali -67 -12024 -34 -11991 0 FreeSerif 160 0 0 0 word169
port 269 nsew
flabel locali -67 -12095 -34 -12062 0 FreeSerif 160 0 0 0 word170
port 270 nsew
flabel locali -67 -12166 -34 -12133 0 FreeSerif 160 0 0 0 word171
port 271 nsew
flabel locali -67 -12237 -34 -12204 0 FreeSerif 160 0 0 0 word172
port 272 nsew
flabel locali -67 -12308 -34 -12275 0 FreeSerif 160 0 0 0 word173
port 273 nsew
flabel locali -67 -12379 -34 -12346 0 FreeSerif 160 0 0 0 word174
port 274 nsew
flabel locali -67 -12450 -34 -12417 0 FreeSerif 160 0 0 0 word175
port 275 nsew
flabel locali -67 -12521 -34 -12488 0 FreeSerif 160 0 0 0 word176
port 276 nsew
flabel locali -67 -12592 -34 -12559 0 FreeSerif 160 0 0 0 word177
port 277 nsew
flabel locali -67 -12663 -34 -12630 0 FreeSerif 160 0 0 0 word178
port 278 nsew
flabel locali -67 -12734 -34 -12701 0 FreeSerif 160 0 0 0 word179
port 279 nsew
flabel locali -67 -12805 -34 -12772 0 FreeSerif 160 0 0 0 word180
port 280 nsew
flabel locali -67 -12876 -34 -12843 0 FreeSerif 160 0 0 0 word181
port 281 nsew
flabel locali -67 -12947 -34 -12914 0 FreeSerif 160 0 0 0 word182
port 282 nsew
flabel locali -67 -13018 -34 -12985 0 FreeSerif 160 0 0 0 word183
port 283 nsew
flabel locali -67 -13089 -34 -13056 0 FreeSerif 160 0 0 0 word184
port 284 nsew
flabel locali -67 -13160 -34 -13127 0 FreeSerif 160 0 0 0 word185
port 285 nsew
flabel locali -67 -13231 -34 -13198 0 FreeSerif 160 0 0 0 word186
port 286 nsew
flabel locali -67 -13302 -34 -13269 0 FreeSerif 160 0 0 0 word187
port 287 nsew
flabel locali -67 -13373 -34 -13340 0 FreeSerif 160 0 0 0 word188
port 288 nsew
flabel locali -67 -13444 -34 -13411 0 FreeSerif 160 0 0 0 word189
port 289 nsew
flabel locali -67 -13515 -34 -13482 0 FreeSerif 160 0 0 0 word190
port 290 nsew
flabel locali -67 -13586 -34 -13553 0 FreeSerif 160 0 0 0 word191
port 291 nsew
flabel locali -67 -13657 -34 -13624 0 FreeSerif 160 0 0 0 word192
port 292 nsew
flabel locali -67 -13728 -34 -13695 0 FreeSerif 160 0 0 0 word193
port 293 nsew
flabel locali -67 -13799 -34 -13766 0 FreeSerif 160 0 0 0 word194
port 294 nsew
flabel locali -67 -13870 -34 -13837 0 FreeSerif 160 0 0 0 word195
port 295 nsew
flabel locali -67 -13941 -34 -13908 0 FreeSerif 160 0 0 0 word196
port 296 nsew
flabel locali -67 -14012 -34 -13979 0 FreeSerif 160 0 0 0 word197
port 297 nsew
flabel locali -67 -14083 -34 -14050 0 FreeSerif 160 0 0 0 word198
port 298 nsew
flabel locali -67 -14154 -34 -14121 0 FreeSerif 160 0 0 0 word199
port 299 nsew
flabel locali -67 -14225 -34 -14192 0 FreeSerif 160 0 0 0 word200
port 300 nsew
flabel locali -67 -14296 -34 -14263 0 FreeSerif 160 0 0 0 word201
port 301 nsew
flabel locali -67 -14367 -34 -14334 0 FreeSerif 160 0 0 0 word202
port 302 nsew
flabel locali -67 -14438 -34 -14405 0 FreeSerif 160 0 0 0 word203
port 303 nsew
flabel locali -67 -14509 -34 -14476 0 FreeSerif 160 0 0 0 word204
port 304 nsew
flabel locali -67 -14580 -34 -14547 0 FreeSerif 160 0 0 0 word205
port 305 nsew
flabel locali -67 -14651 -34 -14618 0 FreeSerif 160 0 0 0 word206
port 306 nsew
flabel locali -67 -14722 -34 -14689 0 FreeSerif 160 0 0 0 word207
port 307 nsew
flabel locali -67 -14793 -34 -14760 0 FreeSerif 160 0 0 0 word208
port 308 nsew
flabel locali -67 -14864 -34 -14831 0 FreeSerif 160 0 0 0 word209
port 309 nsew
flabel locali -67 -14935 -34 -14902 0 FreeSerif 160 0 0 0 word210
port 310 nsew
flabel locali -67 -15006 -34 -14973 0 FreeSerif 160 0 0 0 word211
port 311 nsew
flabel locali -67 -15077 -34 -15044 0 FreeSerif 160 0 0 0 word212
port 312 nsew
flabel locali -67 -15148 -34 -15115 0 FreeSerif 160 0 0 0 word213
port 313 nsew
flabel locali -67 -15219 -34 -15186 0 FreeSerif 160 0 0 0 word214
port 314 nsew
flabel locali -67 -15290 -34 -15257 0 FreeSerif 160 0 0 0 word215
port 315 nsew
flabel locali -67 -15361 -34 -15328 0 FreeSerif 160 0 0 0 word216
port 316 nsew
flabel locali -67 -15432 -34 -15399 0 FreeSerif 160 0 0 0 word217
port 317 nsew
flabel locali -67 -15503 -34 -15470 0 FreeSerif 160 0 0 0 word218
port 318 nsew
flabel locali -67 -15574 -34 -15541 0 FreeSerif 160 0 0 0 word219
port 319 nsew
flabel locali -67 -15645 -34 -15612 0 FreeSerif 160 0 0 0 word220
port 320 nsew
flabel locali -67 -15716 -34 -15683 0 FreeSerif 160 0 0 0 word221
port 321 nsew
flabel locali -67 -15787 -34 -15754 0 FreeSerif 160 0 0 0 word222
port 322 nsew
flabel locali -67 -15858 -34 -15825 0 FreeSerif 160 0 0 0 word223
port 323 nsew
flabel locali -67 -15929 -34 -15896 0 FreeSerif 160 0 0 0 word224
port 324 nsew
flabel locali -67 -16000 -34 -15967 0 FreeSerif 160 0 0 0 word225
port 325 nsew
flabel locali -67 -16071 -34 -16038 0 FreeSerif 160 0 0 0 word226
port 326 nsew
flabel locali -67 -16142 -34 -16109 0 FreeSerif 160 0 0 0 word227
port 327 nsew
flabel locali -67 -16213 -34 -16180 0 FreeSerif 160 0 0 0 word228
port 328 nsew
flabel locali -67 -16284 -34 -16251 0 FreeSerif 160 0 0 0 word229
port 329 nsew
flabel locali -67 -16355 -34 -16322 0 FreeSerif 160 0 0 0 word230
port 330 nsew
flabel locali -67 -16426 -34 -16393 0 FreeSerif 160 0 0 0 word231
port 331 nsew
flabel locali -67 -16497 -34 -16464 0 FreeSerif 160 0 0 0 word232
port 332 nsew
flabel locali -67 -16568 -34 -16535 0 FreeSerif 160 0 0 0 word233
port 333 nsew
flabel locali -67 -16639 -34 -16606 0 FreeSerif 160 0 0 0 word234
port 334 nsew
flabel locali -67 -16710 -34 -16677 0 FreeSerif 160 0 0 0 word235
port 335 nsew
flabel locali -67 -16781 -34 -16748 0 FreeSerif 160 0 0 0 word236
port 336 nsew
flabel locali -67 -16852 -34 -16819 0 FreeSerif 160 0 0 0 word237
port 337 nsew
flabel locali -67 -16923 -34 -16890 0 FreeSerif 160 0 0 0 word238
port 338 nsew
flabel locali -67 -16994 -34 -16961 0 FreeSerif 160 0 0 0 word239
port 339 nsew
flabel locali -67 -17065 -34 -17032 0 FreeSerif 160 0 0 0 word240
port 340 nsew
flabel locali -67 -17136 -34 -17103 0 FreeSerif 160 0 0 0 word241
port 341 nsew
flabel locali -67 -17207 -34 -17174 0 FreeSerif 160 0 0 0 word242
port 342 nsew
flabel locali -67 -17278 -34 -17245 0 FreeSerif 160 0 0 0 word243
port 343 nsew
flabel locali -67 -17349 -34 -17316 0 FreeSerif 160 0 0 0 word244
port 344 nsew
flabel locali -67 -17420 -34 -17387 0 FreeSerif 160 0 0 0 word245
port 345 nsew
flabel locali -67 -17491 -34 -17458 0 FreeSerif 160 0 0 0 word246
port 346 nsew
flabel locali -67 -17562 -34 -17529 0 FreeSerif 160 0 0 0 word247
port 347 nsew
flabel locali -67 -17633 -34 -17600 0 FreeSerif 160 0 0 0 word248
port 348 nsew
flabel locali -67 -17704 -34 -17671 0 FreeSerif 160 0 0 0 word249
port 349 nsew
flabel locali -67 -17775 -34 -17742 0 FreeSerif 160 0 0 0 word250
port 350 nsew
flabel locali -67 -17846 -34 -17813 0 FreeSerif 160 0 0 0 word251
port 351 nsew
flabel locali -67 -17917 -34 -17884 0 FreeSerif 160 0 0 0 word252
port 352 nsew
flabel locali -67 -17988 -34 -17955 0 FreeSerif 160 0 0 0 word253
port 353 nsew
flabel locali -67 -18059 -34 -18026 0 FreeSerif 160 0 0 0 word254
port 354 nsew
flabel locali -67 -18130 -34 -18097 0 FreeSerif 160 0 0 0 word255
port 355 nsew
flabel locali -67 -18201 -34 -18168 0 FreeSerif 160 0 0 0 word256
port 356 nsew
flabel locali -67 -18272 -34 -18239 0 FreeSerif 160 0 0 0 word257
port 357 nsew
flabel locali -67 -18343 -34 -18310 0 FreeSerif 160 0 0 0 word258
port 358 nsew
flabel locali -67 -18414 -34 -18381 0 FreeSerif 160 0 0 0 word259
port 359 nsew
flabel locali -67 -18485 -34 -18452 0 FreeSerif 160 0 0 0 word260
port 360 nsew
flabel locali -67 -18556 -34 -18523 0 FreeSerif 160 0 0 0 word261
port 361 nsew
flabel locali -67 -18627 -34 -18594 0 FreeSerif 160 0 0 0 word262
port 362 nsew
flabel locali -67 -18698 -34 -18665 0 FreeSerif 160 0 0 0 word263
port 363 nsew
flabel locali -67 -18769 -34 -18736 0 FreeSerif 160 0 0 0 word264
port 364 nsew
flabel locali -67 -18840 -34 -18807 0 FreeSerif 160 0 0 0 word265
port 365 nsew
flabel locali -67 -18911 -34 -18878 0 FreeSerif 160 0 0 0 word266
port 366 nsew
flabel locali -67 -18982 -34 -18949 0 FreeSerif 160 0 0 0 word267
port 367 nsew
flabel locali -67 -19053 -34 -19020 0 FreeSerif 160 0 0 0 word268
port 368 nsew
flabel locali -67 -19124 -34 -19091 0 FreeSerif 160 0 0 0 word269
port 369 nsew
flabel locali -67 -19195 -34 -19162 0 FreeSerif 160 0 0 0 word270
port 370 nsew
flabel locali -67 -19266 -34 -19233 0 FreeSerif 160 0 0 0 word271
port 371 nsew
flabel locali -67 -19337 -34 -19304 0 FreeSerif 160 0 0 0 word272
port 372 nsew
flabel locali -67 -19408 -34 -19375 0 FreeSerif 160 0 0 0 word273
port 373 nsew
flabel locali -67 -19479 -34 -19446 0 FreeSerif 160 0 0 0 word274
port 374 nsew
flabel locali -67 -19550 -34 -19517 0 FreeSerif 160 0 0 0 word275
port 375 nsew
flabel locali -67 -19621 -34 -19588 0 FreeSerif 160 0 0 0 word276
port 376 nsew
flabel locali -67 -19692 -34 -19659 0 FreeSerif 160 0 0 0 word277
port 377 nsew
flabel locali -67 -19763 -34 -19730 0 FreeSerif 160 0 0 0 word278
port 378 nsew
flabel locali -67 -19834 -34 -19801 0 FreeSerif 160 0 0 0 word279
port 379 nsew
flabel locali -67 -19905 -34 -19872 0 FreeSerif 160 0 0 0 word280
port 380 nsew
flabel locali -67 -19976 -34 -19943 0 FreeSerif 160 0 0 0 word281
port 381 nsew
flabel locali -67 -20047 -34 -20014 0 FreeSerif 160 0 0 0 word282
port 382 nsew
flabel locali -67 -20118 -34 -20085 0 FreeSerif 160 0 0 0 word283
port 383 nsew
flabel locali -67 -20189 -34 -20156 0 FreeSerif 160 0 0 0 word284
port 384 nsew
flabel locali -67 -20260 -34 -20227 0 FreeSerif 160 0 0 0 word285
port 385 nsew
flabel locali -67 -20331 -34 -20298 0 FreeSerif 160 0 0 0 word286
port 386 nsew
flabel locali -67 -20402 -34 -20369 0 FreeSerif 160 0 0 0 word287
port 387 nsew
flabel locali -67 -20473 -34 -20440 0 FreeSerif 160 0 0 0 word288
port 388 nsew
flabel locali -67 -20544 -34 -20511 0 FreeSerif 160 0 0 0 word289
port 389 nsew
flabel locali -67 -20615 -34 -20582 0 FreeSerif 160 0 0 0 word290
port 390 nsew
flabel locali -67 -20686 -34 -20653 0 FreeSerif 160 0 0 0 word291
port 391 nsew
flabel locali -67 -20757 -34 -20724 0 FreeSerif 160 0 0 0 word292
port 392 nsew
flabel locali -67 -20828 -34 -20795 0 FreeSerif 160 0 0 0 word293
port 393 nsew
flabel locali -67 -20899 -34 -20866 0 FreeSerif 160 0 0 0 word294
port 394 nsew
flabel locali -67 -20970 -34 -20937 0 FreeSerif 160 0 0 0 word295
port 395 nsew
flabel locali -67 -21041 -34 -21008 0 FreeSerif 160 0 0 0 word296
port 396 nsew
flabel locali -67 -21112 -34 -21079 0 FreeSerif 160 0 0 0 word297
port 397 nsew
flabel locali -67 -21183 -34 -21150 0 FreeSerif 160 0 0 0 word298
port 398 nsew
flabel locali -67 -21254 -34 -21221 0 FreeSerif 160 0 0 0 word299
port 399 nsew
flabel locali -67 -21325 -34 -21292 0 FreeSerif 160 0 0 0 word300
port 400 nsew
flabel locali -67 -21396 -34 -21363 0 FreeSerif 160 0 0 0 word301
port 401 nsew
flabel locali -67 -21467 -34 -21434 0 FreeSerif 160 0 0 0 word302
port 402 nsew
flabel locali -67 -21538 -34 -21505 0 FreeSerif 160 0 0 0 word303
port 403 nsew
flabel locali -67 -21609 -34 -21576 0 FreeSerif 160 0 0 0 word304
port 404 nsew
flabel locali -67 -21680 -34 -21647 0 FreeSerif 160 0 0 0 word305
port 405 nsew
flabel locali -67 -21751 -34 -21718 0 FreeSerif 160 0 0 0 word306
port 406 nsew
flabel locali -67 -21822 -34 -21789 0 FreeSerif 160 0 0 0 word307
port 407 nsew
flabel locali -67 -21893 -34 -21860 0 FreeSerif 160 0 0 0 word308
port 408 nsew
flabel locali -67 -21964 -34 -21931 0 FreeSerif 160 0 0 0 word309
port 409 nsew
flabel locali -67 -22035 -34 -22002 0 FreeSerif 160 0 0 0 word310
port 410 nsew
flabel locali -67 -22106 -34 -22073 0 FreeSerif 160 0 0 0 word311
port 411 nsew
flabel locali -67 -22177 -34 -22144 0 FreeSerif 160 0 0 0 word312
port 412 nsew
flabel locali -67 -22248 -34 -22215 0 FreeSerif 160 0 0 0 word313
port 413 nsew
flabel locali -67 -22319 -34 -22286 0 FreeSerif 160 0 0 0 word314
port 414 nsew
flabel locali -67 -22390 -34 -22357 0 FreeSerif 160 0 0 0 word315
port 415 nsew
flabel locali -67 -22461 -34 -22428 0 FreeSerif 160 0 0 0 word316
port 416 nsew
flabel locali -67 -22532 -34 -22499 0 FreeSerif 160 0 0 0 word317
port 417 nsew
flabel locali -67 -22603 -34 -22570 0 FreeSerif 160 0 0 0 word318
port 418 nsew
flabel locali -67 -22674 -34 -22641 0 FreeSerif 160 0 0 0 word319
port 419 nsew
flabel locali -67 -22745 -34 -22712 0 FreeSerif 160 0 0 0 word320
port 420 nsew
flabel locali -67 -22816 -34 -22783 0 FreeSerif 160 0 0 0 word321
port 421 nsew
flabel locali -67 -22887 -34 -22854 0 FreeSerif 160 0 0 0 word322
port 422 nsew
flabel locali -67 -22958 -34 -22925 0 FreeSerif 160 0 0 0 word323
port 423 nsew
flabel locali -67 -23029 -34 -22996 0 FreeSerif 160 0 0 0 word324
port 424 nsew
flabel locali -67 -23100 -34 -23067 0 FreeSerif 160 0 0 0 word325
port 425 nsew
flabel locali -67 -23171 -34 -23138 0 FreeSerif 160 0 0 0 word326
port 426 nsew
flabel locali -67 -23242 -34 -23209 0 FreeSerif 160 0 0 0 word327
port 427 nsew
flabel locali -67 -23313 -34 -23280 0 FreeSerif 160 0 0 0 word328
port 428 nsew
flabel locali -67 -23384 -34 -23351 0 FreeSerif 160 0 0 0 word329
port 429 nsew
flabel locali -67 -23455 -34 -23422 0 FreeSerif 160 0 0 0 word330
port 430 nsew
flabel locali -67 -23526 -34 -23493 0 FreeSerif 160 0 0 0 word331
port 431 nsew
flabel locali -67 -23597 -34 -23564 0 FreeSerif 160 0 0 0 word332
port 432 nsew
flabel locali -67 -23668 -34 -23635 0 FreeSerif 160 0 0 0 word333
port 433 nsew
flabel locali -67 -23739 -34 -23706 0 FreeSerif 160 0 0 0 word334
port 434 nsew
flabel locali -67 -23810 -34 -23777 0 FreeSerif 160 0 0 0 word335
port 435 nsew
flabel locali -67 -23881 -34 -23848 0 FreeSerif 160 0 0 0 word336
port 436 nsew
flabel locali -67 -23952 -34 -23919 0 FreeSerif 160 0 0 0 word337
port 437 nsew
flabel locali -67 -24023 -34 -23990 0 FreeSerif 160 0 0 0 word338
port 438 nsew
flabel locali -67 -24094 -34 -24061 0 FreeSerif 160 0 0 0 word339
port 439 nsew
flabel locali -67 -24165 -34 -24132 0 FreeSerif 160 0 0 0 word340
port 440 nsew
flabel locali -67 -24236 -34 -24203 0 FreeSerif 160 0 0 0 word341
port 441 nsew
flabel locali -67 -24307 -34 -24274 0 FreeSerif 160 0 0 0 word342
port 442 nsew
flabel locali -67 -24378 -34 -24345 0 FreeSerif 160 0 0 0 word343
port 443 nsew
flabel locali -67 -24449 -34 -24416 0 FreeSerif 160 0 0 0 word344
port 444 nsew
flabel locali -67 -24520 -34 -24487 0 FreeSerif 160 0 0 0 word345
port 445 nsew
flabel locali -67 -24591 -34 -24558 0 FreeSerif 160 0 0 0 word346
port 446 nsew
flabel locali -67 -24662 -34 -24629 0 FreeSerif 160 0 0 0 word347
port 447 nsew
flabel locali -67 -24733 -34 -24700 0 FreeSerif 160 0 0 0 word348
port 448 nsew
flabel locali -67 -24804 -34 -24771 0 FreeSerif 160 0 0 0 word349
port 449 nsew
flabel locali -67 -24875 -34 -24842 0 FreeSerif 160 0 0 0 word350
port 450 nsew
flabel locali -67 -24946 -34 -24913 0 FreeSerif 160 0 0 0 word351
port 451 nsew
flabel locali -67 -25017 -34 -24984 0 FreeSerif 160 0 0 0 word352
port 452 nsew
flabel locali -67 -25088 -34 -25055 0 FreeSerif 160 0 0 0 word353
port 453 nsew
flabel locali -67 -25159 -34 -25126 0 FreeSerif 160 0 0 0 word354
port 454 nsew
flabel locali -67 -25230 -34 -25197 0 FreeSerif 160 0 0 0 word355
port 455 nsew
flabel locali -67 -25301 -34 -25268 0 FreeSerif 160 0 0 0 word356
port 456 nsew
flabel locali -67 -25372 -34 -25339 0 FreeSerif 160 0 0 0 word357
port 457 nsew
flabel locali -67 -25443 -34 -25410 0 FreeSerif 160 0 0 0 word358
port 458 nsew
flabel locali -67 -25514 -34 -25481 0 FreeSerif 160 0 0 0 word359
port 459 nsew
flabel locali -67 -25585 -34 -25552 0 FreeSerif 160 0 0 0 word360
port 460 nsew
flabel locali -67 -25656 -34 -25623 0 FreeSerif 160 0 0 0 word361
port 461 nsew
flabel locali -67 -25727 -34 -25694 0 FreeSerif 160 0 0 0 word362
port 462 nsew
flabel locali -67 -25798 -34 -25765 0 FreeSerif 160 0 0 0 word363
port 463 nsew
flabel locali -67 -25869 -34 -25836 0 FreeSerif 160 0 0 0 word364
port 464 nsew
flabel locali -67 -25940 -34 -25907 0 FreeSerif 160 0 0 0 word365
port 465 nsew
flabel locali -67 -26011 -34 -25978 0 FreeSerif 160 0 0 0 word366
port 466 nsew
flabel locali -67 -26082 -34 -26049 0 FreeSerif 160 0 0 0 word367
port 467 nsew
flabel locali -67 -26153 -34 -26120 0 FreeSerif 160 0 0 0 word368
port 468 nsew
flabel locali -67 -26224 -34 -26191 0 FreeSerif 160 0 0 0 word369
port 469 nsew
flabel locali -67 -26295 -34 -26262 0 FreeSerif 160 0 0 0 word370
port 470 nsew
flabel locali -67 -26366 -34 -26333 0 FreeSerif 160 0 0 0 word371
port 471 nsew
flabel locali -67 -26437 -34 -26404 0 FreeSerif 160 0 0 0 word372
port 472 nsew
flabel locali -67 -26508 -34 -26475 0 FreeSerif 160 0 0 0 word373
port 473 nsew
flabel locali -67 -26579 -34 -26546 0 FreeSerif 160 0 0 0 word374
port 474 nsew
flabel locali -67 -26650 -34 -26617 0 FreeSerif 160 0 0 0 word375
port 475 nsew
flabel locali -67 -26721 -34 -26688 0 FreeSerif 160 0 0 0 word376
port 476 nsew
flabel locali -67 -26792 -34 -26759 0 FreeSerif 160 0 0 0 word377
port 477 nsew
flabel locali -67 -26863 -34 -26830 0 FreeSerif 160 0 0 0 word378
port 478 nsew
flabel locali -67 -26934 -34 -26901 0 FreeSerif 160 0 0 0 word379
port 479 nsew
flabel locali -67 -27005 -34 -26972 0 FreeSerif 160 0 0 0 word380
port 480 nsew
flabel locali -67 -27076 -34 -27043 0 FreeSerif 160 0 0 0 word381
port 481 nsew
flabel locali -67 -27147 -34 -27114 0 FreeSerif 160 0 0 0 word382
port 482 nsew
flabel locali -67 -27218 -34 -27185 0 FreeSerif 160 0 0 0 word383
port 483 nsew
flabel locali -67 -27289 -34 -27256 0 FreeSerif 160 0 0 0 word384
port 484 nsew
flabel locali -67 -27360 -34 -27327 0 FreeSerif 160 0 0 0 word385
port 485 nsew
flabel locali -67 -27431 -34 -27398 0 FreeSerif 160 0 0 0 word386
port 486 nsew
flabel locali -67 -27502 -34 -27469 0 FreeSerif 160 0 0 0 word387
port 487 nsew
flabel locali -67 -27573 -34 -27540 0 FreeSerif 160 0 0 0 word388
port 488 nsew
flabel locali -67 -27644 -34 -27611 0 FreeSerif 160 0 0 0 word389
port 489 nsew
flabel locali -67 -27715 -34 -27682 0 FreeSerif 160 0 0 0 word390
port 490 nsew
flabel locali -67 -27786 -34 -27753 0 FreeSerif 160 0 0 0 word391
port 491 nsew
flabel locali -67 -27857 -34 -27824 0 FreeSerif 160 0 0 0 word392
port 492 nsew
flabel locali -67 -27928 -34 -27895 0 FreeSerif 160 0 0 0 word393
port 493 nsew
flabel locali -67 -27999 -34 -27966 0 FreeSerif 160 0 0 0 word394
port 494 nsew
flabel locali -67 -28070 -34 -28037 0 FreeSerif 160 0 0 0 word395
port 495 nsew
flabel locali -67 -28141 -34 -28108 0 FreeSerif 160 0 0 0 word396
port 496 nsew
flabel locali -67 -28212 -34 -28179 0 FreeSerif 160 0 0 0 word397
port 497 nsew
flabel locali -67 -28283 -34 -28250 0 FreeSerif 160 0 0 0 word398
port 498 nsew
flabel locali -67 -28354 -34 -28321 0 FreeSerif 160 0 0 0 word399
port 499 nsew
flabel locali -67 -28425 -34 -28392 0 FreeSerif 160 0 0 0 word400
port 500 nsew
flabel locali -67 -28496 -34 -28463 0 FreeSerif 160 0 0 0 word401
port 501 nsew
flabel locali -67 -28567 -34 -28534 0 FreeSerif 160 0 0 0 word402
port 502 nsew
flabel locali -67 -28638 -34 -28605 0 FreeSerif 160 0 0 0 word403
port 503 nsew
flabel locali -67 -28709 -34 -28676 0 FreeSerif 160 0 0 0 word404
port 504 nsew
flabel locali -67 -28780 -34 -28747 0 FreeSerif 160 0 0 0 word405
port 505 nsew
flabel locali -67 -28851 -34 -28818 0 FreeSerif 160 0 0 0 word406
port 506 nsew
flabel locali -67 -28922 -34 -28889 0 FreeSerif 160 0 0 0 word407
port 507 nsew
flabel locali -67 -28993 -34 -28960 0 FreeSerif 160 0 0 0 word408
port 508 nsew
flabel locali -67 -29064 -34 -29031 0 FreeSerif 160 0 0 0 word409
port 509 nsew
flabel locali -67 -29135 -34 -29102 0 FreeSerif 160 0 0 0 word410
port 510 nsew
flabel locali -67 -29206 -34 -29173 0 FreeSerif 160 0 0 0 word411
port 511 nsew
flabel locali -67 -29277 -34 -29244 0 FreeSerif 160 0 0 0 word412
port 512 nsew
flabel locali -67 -29348 -34 -29315 0 FreeSerif 160 0 0 0 word413
port 513 nsew
flabel locali -67 -29419 -34 -29386 0 FreeSerif 160 0 0 0 word414
port 514 nsew
flabel locali -67 -29490 -34 -29457 0 FreeSerif 160 0 0 0 word415
port 515 nsew
flabel locali -67 -29561 -34 -29528 0 FreeSerif 160 0 0 0 word416
port 516 nsew
flabel locali -67 -29632 -34 -29599 0 FreeSerif 160 0 0 0 word417
port 517 nsew
flabel locali -67 -29703 -34 -29670 0 FreeSerif 160 0 0 0 word418
port 518 nsew
flabel locali -67 -29774 -34 -29741 0 FreeSerif 160 0 0 0 word419
port 519 nsew
flabel locali -67 -29845 -34 -29812 0 FreeSerif 160 0 0 0 word420
port 520 nsew
flabel locali -67 -29916 -34 -29883 0 FreeSerif 160 0 0 0 word421
port 521 nsew
flabel locali -67 -29987 -34 -29954 0 FreeSerif 160 0 0 0 word422
port 522 nsew
flabel locali -67 -30058 -34 -30025 0 FreeSerif 160 0 0 0 word423
port 523 nsew
flabel locali -67 -30129 -34 -30096 0 FreeSerif 160 0 0 0 word424
port 524 nsew
flabel locali -67 -30200 -34 -30167 0 FreeSerif 160 0 0 0 word425
port 525 nsew
flabel locali -67 -30271 -34 -30238 0 FreeSerif 160 0 0 0 word426
port 526 nsew
flabel locali -67 -30342 -34 -30309 0 FreeSerif 160 0 0 0 word427
port 527 nsew
flabel locali -67 -30413 -34 -30380 0 FreeSerif 160 0 0 0 word428
port 528 nsew
flabel locali -67 -30484 -34 -30451 0 FreeSerif 160 0 0 0 word429
port 529 nsew
flabel locali -67 -30555 -34 -30522 0 FreeSerif 160 0 0 0 word430
port 530 nsew
flabel locali -67 -30626 -34 -30593 0 FreeSerif 160 0 0 0 word431
port 531 nsew
flabel locali -67 -30697 -34 -30664 0 FreeSerif 160 0 0 0 word432
port 532 nsew
flabel locali -67 -30768 -34 -30735 0 FreeSerif 160 0 0 0 word433
port 533 nsew
flabel locali -67 -30839 -34 -30806 0 FreeSerif 160 0 0 0 word434
port 534 nsew
flabel locali -67 -30910 -34 -30877 0 FreeSerif 160 0 0 0 word435
port 535 nsew
flabel locali -67 -30981 -34 -30948 0 FreeSerif 160 0 0 0 word436
port 536 nsew
flabel locali -67 -31052 -34 -31019 0 FreeSerif 160 0 0 0 word437
port 537 nsew
flabel locali -67 -31123 -34 -31090 0 FreeSerif 160 0 0 0 word438
port 538 nsew
flabel locali -67 -31194 -34 -31161 0 FreeSerif 160 0 0 0 word439
port 539 nsew
flabel locali -67 -31265 -34 -31232 0 FreeSerif 160 0 0 0 word440
port 540 nsew
flabel locali -67 -31336 -34 -31303 0 FreeSerif 160 0 0 0 word441
port 541 nsew
flabel locali -67 -31407 -34 -31374 0 FreeSerif 160 0 0 0 word442
port 542 nsew
flabel locali -67 -31478 -34 -31445 0 FreeSerif 160 0 0 0 word443
port 543 nsew
flabel locali -67 -31549 -34 -31516 0 FreeSerif 160 0 0 0 word444
port 544 nsew
flabel locali -67 -31620 -34 -31587 0 FreeSerif 160 0 0 0 word445
port 545 nsew
flabel locali -67 -31691 -34 -31658 0 FreeSerif 160 0 0 0 word446
port 546 nsew
flabel locali -67 -31762 -34 -31729 0 FreeSerif 160 0 0 0 word447
port 547 nsew
flabel locali -67 -31833 -34 -31800 0 FreeSerif 160 0 0 0 word448
port 548 nsew
flabel locali -67 -31904 -34 -31871 0 FreeSerif 160 0 0 0 word449
port 549 nsew
flabel locali -67 -31975 -34 -31942 0 FreeSerif 160 0 0 0 word450
port 550 nsew
flabel locali -67 -32046 -34 -32013 0 FreeSerif 160 0 0 0 word451
port 551 nsew
flabel locali -67 -32117 -34 -32084 0 FreeSerif 160 0 0 0 word452
port 552 nsew
flabel locali -67 -32188 -34 -32155 0 FreeSerif 160 0 0 0 word453
port 553 nsew
flabel locali -67 -32259 -34 -32226 0 FreeSerif 160 0 0 0 word454
port 554 nsew
flabel locali -67 -32330 -34 -32297 0 FreeSerif 160 0 0 0 word455
port 555 nsew
flabel locali -67 -32401 -34 -32368 0 FreeSerif 160 0 0 0 word456
port 556 nsew
flabel locali -67 -32472 -34 -32439 0 FreeSerif 160 0 0 0 word457
port 557 nsew
flabel locali -67 -32543 -34 -32510 0 FreeSerif 160 0 0 0 word458
port 558 nsew
flabel locali -67 -32614 -34 -32581 0 FreeSerif 160 0 0 0 word459
port 559 nsew
flabel locali -67 -32685 -34 -32652 0 FreeSerif 160 0 0 0 word460
port 560 nsew
flabel locali -67 -32756 -34 -32723 0 FreeSerif 160 0 0 0 word461
port 561 nsew
flabel locali -67 -32827 -34 -32794 0 FreeSerif 160 0 0 0 word462
port 562 nsew
flabel locali -67 -32898 -34 -32865 0 FreeSerif 160 0 0 0 word463
port 563 nsew
flabel locali -67 -32969 -34 -32936 0 FreeSerif 160 0 0 0 word464
port 564 nsew
flabel locali -67 -33040 -34 -33007 0 FreeSerif 160 0 0 0 word465
port 565 nsew
flabel locali -67 -33111 -34 -33078 0 FreeSerif 160 0 0 0 word466
port 566 nsew
flabel locali -67 -33182 -34 -33149 0 FreeSerif 160 0 0 0 word467
port 567 nsew
flabel locali -67 -33253 -34 -33220 0 FreeSerif 160 0 0 0 word468
port 568 nsew
flabel locali -67 -33324 -34 -33291 0 FreeSerif 160 0 0 0 word469
port 569 nsew
flabel locali -67 -33395 -34 -33362 0 FreeSerif 160 0 0 0 word470
port 570 nsew
flabel locali -67 -33466 -34 -33433 0 FreeSerif 160 0 0 0 word471
port 571 nsew
flabel locali -67 -33537 -34 -33504 0 FreeSerif 160 0 0 0 word472
port 572 nsew
flabel locali -67 -33608 -34 -33575 0 FreeSerif 160 0 0 0 word473
port 573 nsew
flabel locali -67 -33679 -34 -33646 0 FreeSerif 160 0 0 0 word474
port 574 nsew
flabel locali -67 -33750 -34 -33717 0 FreeSerif 160 0 0 0 word475
port 575 nsew
flabel locali -67 -33821 -34 -33788 0 FreeSerif 160 0 0 0 word476
port 576 nsew
flabel locali -67 -33892 -34 -33859 0 FreeSerif 160 0 0 0 word477
port 577 nsew
flabel locali -67 -33963 -34 -33930 0 FreeSerif 160 0 0 0 word478
port 578 nsew
flabel locali -67 -34034 -34 -34001 0 FreeSerif 160 0 0 0 word479
port 579 nsew
flabel locali -67 -34105 -34 -34072 0 FreeSerif 160 0 0 0 word480
port 580 nsew
flabel locali -67 -34176 -34 -34143 0 FreeSerif 160 0 0 0 word481
port 581 nsew
flabel locali -67 -34247 -34 -34214 0 FreeSerif 160 0 0 0 word482
port 582 nsew
flabel locali -67 -34318 -34 -34285 0 FreeSerif 160 0 0 0 word483
port 583 nsew
flabel locali -67 -34389 -34 -34356 0 FreeSerif 160 0 0 0 word484
port 584 nsew
flabel locali -67 -34460 -34 -34427 0 FreeSerif 160 0 0 0 word485
port 585 nsew
flabel locali -67 -34531 -34 -34498 0 FreeSerif 160 0 0 0 word486
port 586 nsew
flabel locali -67 -34602 -34 -34569 0 FreeSerif 160 0 0 0 word487
port 587 nsew
flabel locali -67 -34673 -34 -34640 0 FreeSerif 160 0 0 0 word488
port 588 nsew
flabel locali -67 -34744 -34 -34711 0 FreeSerif 160 0 0 0 word489
port 589 nsew
flabel locali -67 -34815 -34 -34782 0 FreeSerif 160 0 0 0 word490
port 590 nsew
flabel locali -67 -34886 -34 -34853 0 FreeSerif 160 0 0 0 word491
port 591 nsew
flabel locali -67 -34957 -34 -34924 0 FreeSerif 160 0 0 0 word492
port 592 nsew
flabel locali -67 -35028 -34 -34995 0 FreeSerif 160 0 0 0 word493
port 593 nsew
flabel locali -67 -35099 -34 -35066 0 FreeSerif 160 0 0 0 word494
port 594 nsew
flabel locali -67 -35170 -34 -35137 0 FreeSerif 160 0 0 0 word495
port 595 nsew
flabel locali -67 -35241 -34 -35208 0 FreeSerif 160 0 0 0 word496
port 596 nsew
flabel locali -67 -35312 -34 -35279 0 FreeSerif 160 0 0 0 word497
port 597 nsew
flabel locali -67 -35383 -34 -35350 0 FreeSerif 160 0 0 0 word498
port 598 nsew
flabel locali -67 -35454 -34 -35421 0 FreeSerif 160 0 0 0 word499
port 599 nsew
flabel locali -67 -35525 -34 -35492 0 FreeSerif 160 0 0 0 word500
port 600 nsew
flabel locali -67 -35596 -34 -35563 0 FreeSerif 160 0 0 0 word501
port 601 nsew
flabel locali -67 -35667 -34 -35634 0 FreeSerif 160 0 0 0 word502
port 602 nsew
flabel locali -67 -35738 -34 -35705 0 FreeSerif 160 0 0 0 word503
port 603 nsew
flabel locali -67 -35809 -34 -35776 0 FreeSerif 160 0 0 0 word504
port 604 nsew
flabel locali -67 -35880 -34 -35847 0 FreeSerif 160 0 0 0 word505
port 605 nsew
flabel locali -67 -35951 -34 -35918 0 FreeSerif 160 0 0 0 word506
port 606 nsew
flabel locali -67 -36022 -34 -35989 0 FreeSerif 160 0 0 0 word507
port 607 nsew
flabel locali -67 -36093 -34 -36060 0 FreeSerif 160 0 0 0 word508
port 608 nsew
flabel locali -67 -36164 -34 -36131 0 FreeSerif 160 0 0 0 word509
port 609 nsew
flabel locali -67 -36235 -34 -36202 0 FreeSerif 160 0 0 0 word510
port 610 nsew
flabel locali -67 -36306 -34 -36273 0 FreeSerif 160 0 0 0 word511
port 611 nsew
flabel locali -67 -36377 -34 -36344 0 FreeSerif 160 0 0 0 word512
port 612 nsew
flabel locali -67 -36448 -34 -36415 0 FreeSerif 160 0 0 0 word513
port 613 nsew
flabel locali -67 -36519 -34 -36486 0 FreeSerif 160 0 0 0 word514
port 614 nsew
flabel locali -67 -36590 -34 -36557 0 FreeSerif 160 0 0 0 word515
port 615 nsew
flabel locali -67 -36661 -34 -36628 0 FreeSerif 160 0 0 0 word516
port 616 nsew
flabel locali -67 -36732 -34 -36699 0 FreeSerif 160 0 0 0 word517
port 617 nsew
flabel locali -67 -36803 -34 -36770 0 FreeSerif 160 0 0 0 word518
port 618 nsew
flabel locali -67 -36874 -34 -36841 0 FreeSerif 160 0 0 0 word519
port 619 nsew
flabel locali -67 -36945 -34 -36912 0 FreeSerif 160 0 0 0 word520
port 620 nsew
flabel locali -67 -37016 -34 -36983 0 FreeSerif 160 0 0 0 word521
port 621 nsew
flabel locali -67 -37087 -34 -37054 0 FreeSerif 160 0 0 0 word522
port 622 nsew
flabel locali -67 -37158 -34 -37125 0 FreeSerif 160 0 0 0 word523
port 623 nsew
flabel locali -67 -37229 -34 -37196 0 FreeSerif 160 0 0 0 word524
port 624 nsew
flabel locali -67 -37300 -34 -37267 0 FreeSerif 160 0 0 0 word525
port 625 nsew
flabel locali -67 -37371 -34 -37338 0 FreeSerif 160 0 0 0 word526
port 626 nsew
flabel locali -67 -37442 -34 -37409 0 FreeSerif 160 0 0 0 word527
port 627 nsew
flabel locali -67 -37513 -34 -37480 0 FreeSerif 160 0 0 0 word528
port 628 nsew
flabel locali -67 -37584 -34 -37551 0 FreeSerif 160 0 0 0 word529
port 629 nsew
flabel locali -67 -37655 -34 -37622 0 FreeSerif 160 0 0 0 word530
port 630 nsew
flabel locali -67 -37726 -34 -37693 0 FreeSerif 160 0 0 0 word531
port 631 nsew
flabel locali -67 -37797 -34 -37764 0 FreeSerif 160 0 0 0 word532
port 632 nsew
flabel locali -67 -37868 -34 -37835 0 FreeSerif 160 0 0 0 word533
port 633 nsew
flabel locali -67 -37939 -34 -37906 0 FreeSerif 160 0 0 0 word534
port 634 nsew
flabel locali -67 -38010 -34 -37977 0 FreeSerif 160 0 0 0 word535
port 635 nsew
flabel locali -67 -38081 -34 -38048 0 FreeSerif 160 0 0 0 word536
port 636 nsew
flabel locali -67 -38152 -34 -38119 0 FreeSerif 160 0 0 0 word537
port 637 nsew
flabel locali -67 -38223 -34 -38190 0 FreeSerif 160 0 0 0 word538
port 638 nsew
flabel locali -67 -38294 -34 -38261 0 FreeSerif 160 0 0 0 word539
port 639 nsew
flabel locali -67 -38365 -34 -38332 0 FreeSerif 160 0 0 0 word540
port 640 nsew
flabel locali -67 -38436 -34 -38403 0 FreeSerif 160 0 0 0 word541
port 641 nsew
flabel locali -67 -38507 -34 -38474 0 FreeSerif 160 0 0 0 word542
port 642 nsew
flabel locali -67 -38578 -34 -38545 0 FreeSerif 160 0 0 0 word543
port 643 nsew
flabel locali -67 -38649 -34 -38616 0 FreeSerif 160 0 0 0 word544
port 644 nsew
flabel locali -67 -38720 -34 -38687 0 FreeSerif 160 0 0 0 word545
port 645 nsew
flabel locali -67 -38791 -34 -38758 0 FreeSerif 160 0 0 0 word546
port 646 nsew
flabel locali -67 -38862 -34 -38829 0 FreeSerif 160 0 0 0 word547
port 647 nsew
flabel locali -67 -38933 -34 -38900 0 FreeSerif 160 0 0 0 word548
port 648 nsew
flabel locali -67 -39004 -34 -38971 0 FreeSerif 160 0 0 0 word549
port 649 nsew
flabel locali -67 -39075 -34 -39042 0 FreeSerif 160 0 0 0 word550
port 650 nsew
flabel locali -67 -39146 -34 -39113 0 FreeSerif 160 0 0 0 word551
port 651 nsew
flabel locali -67 -39217 -34 -39184 0 FreeSerif 160 0 0 0 word552
port 652 nsew
flabel locali -67 -39288 -34 -39255 0 FreeSerif 160 0 0 0 word553
port 653 nsew
flabel locali -67 -39359 -34 -39326 0 FreeSerif 160 0 0 0 word554
port 654 nsew
flabel locali -67 -39430 -34 -39397 0 FreeSerif 160 0 0 0 word555
port 655 nsew
flabel locali -67 -39501 -34 -39468 0 FreeSerif 160 0 0 0 word556
port 656 nsew
flabel locali -67 -39572 -34 -39539 0 FreeSerif 160 0 0 0 word557
port 657 nsew
flabel locali -67 -39643 -34 -39610 0 FreeSerif 160 0 0 0 word558
port 658 nsew
flabel locali -67 -39714 -34 -39681 0 FreeSerif 160 0 0 0 word559
port 659 nsew
flabel locali -67 -39785 -34 -39752 0 FreeSerif 160 0 0 0 word560
port 660 nsew
flabel locali -67 -39856 -34 -39823 0 FreeSerif 160 0 0 0 word561
port 661 nsew
flabel locali -67 -39927 -34 -39894 0 FreeSerif 160 0 0 0 word562
port 662 nsew
flabel locali -67 -39998 -34 -39965 0 FreeSerif 160 0 0 0 word563
port 663 nsew
flabel locali -67 -40069 -34 -40036 0 FreeSerif 160 0 0 0 word564
port 664 nsew
flabel locali -67 -40140 -34 -40107 0 FreeSerif 160 0 0 0 word565
port 665 nsew
flabel locali -67 -40211 -34 -40178 0 FreeSerif 160 0 0 0 word566
port 666 nsew
flabel locali -67 -40282 -34 -40249 0 FreeSerif 160 0 0 0 word567
port 667 nsew
flabel locali -67 -40353 -34 -40320 0 FreeSerif 160 0 0 0 word568
port 668 nsew
flabel locali -67 -40424 -34 -40391 0 FreeSerif 160 0 0 0 word569
port 669 nsew
flabel locali -67 -40495 -34 -40462 0 FreeSerif 160 0 0 0 word570
port 670 nsew
flabel locali -67 -40566 -34 -40533 0 FreeSerif 160 0 0 0 word571
port 671 nsew
flabel locali -67 -40637 -34 -40604 0 FreeSerif 160 0 0 0 word572
port 672 nsew
flabel locali -67 -40708 -34 -40675 0 FreeSerif 160 0 0 0 word573
port 673 nsew
flabel locali -67 -40779 -34 -40746 0 FreeSerif 160 0 0 0 word574
port 674 nsew
flabel locali -67 -40850 -34 -40817 0 FreeSerif 160 0 0 0 word575
port 675 nsew
flabel locali -67 -40921 -34 -40888 0 FreeSerif 160 0 0 0 word576
port 676 nsew
flabel locali -67 -40992 -34 -40959 0 FreeSerif 160 0 0 0 word577
port 677 nsew
flabel locali -67 -41063 -34 -41030 0 FreeSerif 160 0 0 0 word578
port 678 nsew
flabel locali -67 -41134 -34 -41101 0 FreeSerif 160 0 0 0 word579
port 679 nsew
flabel locali -67 -41205 -34 -41172 0 FreeSerif 160 0 0 0 word580
port 680 nsew
flabel locali -67 -41276 -34 -41243 0 FreeSerif 160 0 0 0 word581
port 681 nsew
flabel locali -67 -41347 -34 -41314 0 FreeSerif 160 0 0 0 word582
port 682 nsew
flabel locali -67 -41418 -34 -41385 0 FreeSerif 160 0 0 0 word583
port 683 nsew
flabel locali -67 -41489 -34 -41456 0 FreeSerif 160 0 0 0 word584
port 684 nsew
flabel locali -67 -41560 -34 -41527 0 FreeSerif 160 0 0 0 word585
port 685 nsew
flabel locali -67 -41631 -34 -41598 0 FreeSerif 160 0 0 0 word586
port 686 nsew
flabel locali -67 -41702 -34 -41669 0 FreeSerif 160 0 0 0 word587
port 687 nsew
flabel locali -67 -41773 -34 -41740 0 FreeSerif 160 0 0 0 word588
port 688 nsew
flabel locali -67 -41844 -34 -41811 0 FreeSerif 160 0 0 0 word589
port 689 nsew
flabel locali -67 -41915 -34 -41882 0 FreeSerif 160 0 0 0 word590
port 690 nsew
flabel locali -67 -41986 -34 -41953 0 FreeSerif 160 0 0 0 word591
port 691 nsew
flabel locali -67 -42057 -34 -42024 0 FreeSerif 160 0 0 0 word592
port 692 nsew
flabel locali -67 -42128 -34 -42095 0 FreeSerif 160 0 0 0 word593
port 693 nsew
flabel locali -67 -42199 -34 -42166 0 FreeSerif 160 0 0 0 word594
port 694 nsew
flabel locali -67 -42270 -34 -42237 0 FreeSerif 160 0 0 0 word595
port 695 nsew
flabel locali -67 -42341 -34 -42308 0 FreeSerif 160 0 0 0 word596
port 696 nsew
flabel locali -67 -42412 -34 -42379 0 FreeSerif 160 0 0 0 word597
port 697 nsew
flabel locali -67 -42483 -34 -42450 0 FreeSerif 160 0 0 0 word598
port 698 nsew
flabel locali -67 -42554 -34 -42521 0 FreeSerif 160 0 0 0 word599
port 699 nsew
flabel locali -67 -42625 -34 -42592 0 FreeSerif 160 0 0 0 word600
port 700 nsew
flabel locali -67 -42696 -34 -42663 0 FreeSerif 160 0 0 0 word601
port 701 nsew
flabel locali -67 -42767 -34 -42734 0 FreeSerif 160 0 0 0 word602
port 702 nsew
flabel locali -67 -42838 -34 -42805 0 FreeSerif 160 0 0 0 word603
port 703 nsew
flabel locali -67 -42909 -34 -42876 0 FreeSerif 160 0 0 0 word604
port 704 nsew
flabel locali -67 -42980 -34 -42947 0 FreeSerif 160 0 0 0 word605
port 705 nsew
flabel locali -67 -43051 -34 -43018 0 FreeSerif 160 0 0 0 word606
port 706 nsew
flabel locali -67 -43122 -34 -43089 0 FreeSerif 160 0 0 0 word607
port 707 nsew
flabel locali -67 -43193 -34 -43160 0 FreeSerif 160 0 0 0 word608
port 708 nsew
flabel locali -67 -43264 -34 -43231 0 FreeSerif 160 0 0 0 word609
port 709 nsew
flabel locali -67 -43335 -34 -43302 0 FreeSerif 160 0 0 0 word610
port 710 nsew
flabel locali -67 -43406 -34 -43373 0 FreeSerif 160 0 0 0 word611
port 711 nsew
flabel locali -67 -43477 -34 -43444 0 FreeSerif 160 0 0 0 word612
port 712 nsew
flabel locali -67 -43548 -34 -43515 0 FreeSerif 160 0 0 0 word613
port 713 nsew
flabel locali -67 -43619 -34 -43586 0 FreeSerif 160 0 0 0 word614
port 714 nsew
flabel locali -67 -43690 -34 -43657 0 FreeSerif 160 0 0 0 word615
port 715 nsew
flabel locali -67 -43761 -34 -43728 0 FreeSerif 160 0 0 0 word616
port 716 nsew
flabel locali -67 -43832 -34 -43799 0 FreeSerif 160 0 0 0 word617
port 717 nsew
flabel locali -67 -43903 -34 -43870 0 FreeSerif 160 0 0 0 word618
port 718 nsew
flabel locali -67 -43974 -34 -43941 0 FreeSerif 160 0 0 0 word619
port 719 nsew
flabel locali -67 -44045 -34 -44012 0 FreeSerif 160 0 0 0 word620
port 720 nsew
flabel locali -67 -44116 -34 -44083 0 FreeSerif 160 0 0 0 word621
port 721 nsew
flabel locali -67 -44187 -34 -44154 0 FreeSerif 160 0 0 0 word622
port 722 nsew
flabel locali -67 -44258 -34 -44225 0 FreeSerif 160 0 0 0 word623
port 723 nsew
flabel locali -67 -44329 -34 -44296 0 FreeSerif 160 0 0 0 word624
port 724 nsew
flabel locali -67 -44400 -34 -44367 0 FreeSerif 160 0 0 0 word625
port 725 nsew
flabel locali -67 -44471 -34 -44438 0 FreeSerif 160 0 0 0 word626
port 726 nsew
flabel locali -67 -44542 -34 -44509 0 FreeSerif 160 0 0 0 word627
port 727 nsew
flabel locali -67 -44613 -34 -44580 0 FreeSerif 160 0 0 0 word628
port 728 nsew
flabel locali -67 -44684 -34 -44651 0 FreeSerif 160 0 0 0 word629
port 729 nsew
flabel locali -67 -44755 -34 -44722 0 FreeSerif 160 0 0 0 word630
port 730 nsew
flabel locali -67 -44826 -34 -44793 0 FreeSerif 160 0 0 0 word631
port 731 nsew
flabel locali -67 -44897 -34 -44864 0 FreeSerif 160 0 0 0 word632
port 732 nsew
flabel locali -67 -44968 -34 -44935 0 FreeSerif 160 0 0 0 word633
port 733 nsew
flabel locali -67 -45039 -34 -45006 0 FreeSerif 160 0 0 0 word634
port 734 nsew
flabel locali -67 -45110 -34 -45077 0 FreeSerif 160 0 0 0 word635
port 735 nsew
flabel locali -67 -45181 -34 -45148 0 FreeSerif 160 0 0 0 word636
port 736 nsew
flabel locali -67 -45252 -34 -45219 0 FreeSerif 160 0 0 0 word637
port 737 nsew
flabel locali -67 -45323 -34 -45290 0 FreeSerif 160 0 0 0 word638
port 738 nsew
flabel locali -67 -45394 -34 -45361 0 FreeSerif 160 0 0 0 word639
port 739 nsew
flabel locali -67 -45465 -34 -45432 0 FreeSerif 160 0 0 0 word640
port 740 nsew
flabel locali -67 -45536 -34 -45503 0 FreeSerif 160 0 0 0 word641
port 741 nsew
flabel locali -67 -45607 -34 -45574 0 FreeSerif 160 0 0 0 word642
port 742 nsew
flabel locali -67 -45678 -34 -45645 0 FreeSerif 160 0 0 0 word643
port 743 nsew
flabel locali -67 -45749 -34 -45716 0 FreeSerif 160 0 0 0 word644
port 744 nsew
flabel locali -67 -45820 -34 -45787 0 FreeSerif 160 0 0 0 word645
port 745 nsew
flabel locali -67 -45891 -34 -45858 0 FreeSerif 160 0 0 0 word646
port 746 nsew
flabel locali -67 -45962 -34 -45929 0 FreeSerif 160 0 0 0 word647
port 747 nsew
flabel locali -67 -46033 -34 -46000 0 FreeSerif 160 0 0 0 word648
port 748 nsew
flabel locali -67 -46104 -34 -46071 0 FreeSerif 160 0 0 0 word649
port 749 nsew
flabel locali -67 -46175 -34 -46142 0 FreeSerif 160 0 0 0 word650
port 750 nsew
flabel locali -67 -46246 -34 -46213 0 FreeSerif 160 0 0 0 word651
port 751 nsew
flabel locali -67 -46317 -34 -46284 0 FreeSerif 160 0 0 0 word652
port 752 nsew
flabel locali -67 -46388 -34 -46355 0 FreeSerif 160 0 0 0 word653
port 753 nsew
flabel locali -67 -46459 -34 -46426 0 FreeSerif 160 0 0 0 word654
port 754 nsew
flabel locali -67 -46530 -34 -46497 0 FreeSerif 160 0 0 0 word655
port 755 nsew
flabel locali -67 -46601 -34 -46568 0 FreeSerif 160 0 0 0 word656
port 756 nsew
flabel locali -67 -46672 -34 -46639 0 FreeSerif 160 0 0 0 word657
port 757 nsew
flabel locali -67 -46743 -34 -46710 0 FreeSerif 160 0 0 0 word658
port 758 nsew
flabel locali -67 -46814 -34 -46781 0 FreeSerif 160 0 0 0 word659
port 759 nsew
flabel locali -67 -46885 -34 -46852 0 FreeSerif 160 0 0 0 word660
port 760 nsew
flabel locali -67 -46956 -34 -46923 0 FreeSerif 160 0 0 0 word661
port 761 nsew
flabel locali -67 -47027 -34 -46994 0 FreeSerif 160 0 0 0 word662
port 762 nsew
flabel locali -67 -47098 -34 -47065 0 FreeSerif 160 0 0 0 word663
port 763 nsew
flabel locali -67 -47169 -34 -47136 0 FreeSerif 160 0 0 0 word664
port 764 nsew
flabel locali -67 -47240 -34 -47207 0 FreeSerif 160 0 0 0 word665
port 765 nsew
flabel locali -67 -47311 -34 -47278 0 FreeSerif 160 0 0 0 word666
port 766 nsew
flabel locali -67 -47382 -34 -47349 0 FreeSerif 160 0 0 0 word667
port 767 nsew
flabel locali -67 -47453 -34 -47420 0 FreeSerif 160 0 0 0 word668
port 768 nsew
flabel locali -67 -47524 -34 -47491 0 FreeSerif 160 0 0 0 word669
port 769 nsew
flabel locali -67 -47595 -34 -47562 0 FreeSerif 160 0 0 0 word670
port 770 nsew
flabel locali -67 -47666 -34 -47633 0 FreeSerif 160 0 0 0 word671
port 771 nsew
flabel locali -67 -47737 -34 -47704 0 FreeSerif 160 0 0 0 word672
port 772 nsew
flabel locali -67 -47808 -34 -47775 0 FreeSerif 160 0 0 0 word673
port 773 nsew
flabel locali -67 -47879 -34 -47846 0 FreeSerif 160 0 0 0 word674
port 774 nsew
flabel locali -67 -47950 -34 -47917 0 FreeSerif 160 0 0 0 word675
port 775 nsew
flabel locali -67 -48021 -34 -47988 0 FreeSerif 160 0 0 0 word676
port 776 nsew
flabel locali -67 -48092 -34 -48059 0 FreeSerif 160 0 0 0 word677
port 777 nsew
flabel locali -67 -48163 -34 -48130 0 FreeSerif 160 0 0 0 word678
port 778 nsew
flabel locali -67 -48234 -34 -48201 0 FreeSerif 160 0 0 0 word679
port 779 nsew
flabel locali -67 -48305 -34 -48272 0 FreeSerif 160 0 0 0 word680
port 780 nsew
flabel locali -67 -48376 -34 -48343 0 FreeSerif 160 0 0 0 word681
port 781 nsew
flabel locali -67 -48447 -34 -48414 0 FreeSerif 160 0 0 0 word682
port 782 nsew
flabel locali -67 -48518 -34 -48485 0 FreeSerif 160 0 0 0 word683
port 783 nsew
flabel locali -67 -48589 -34 -48556 0 FreeSerif 160 0 0 0 word684
port 784 nsew
flabel locali -67 -48660 -34 -48627 0 FreeSerif 160 0 0 0 word685
port 785 nsew
flabel locali -67 -48731 -34 -48698 0 FreeSerif 160 0 0 0 word686
port 786 nsew
flabel locali -67 -48802 -34 -48769 0 FreeSerif 160 0 0 0 word687
port 787 nsew
flabel locali -67 -48873 -34 -48840 0 FreeSerif 160 0 0 0 word688
port 788 nsew
flabel locali -67 -48944 -34 -48911 0 FreeSerif 160 0 0 0 word689
port 789 nsew
flabel locali -67 -49015 -34 -48982 0 FreeSerif 160 0 0 0 word690
port 790 nsew
flabel locali -67 -49086 -34 -49053 0 FreeSerif 160 0 0 0 word691
port 791 nsew
flabel locali -67 -49157 -34 -49124 0 FreeSerif 160 0 0 0 word692
port 792 nsew
flabel locali -67 -49228 -34 -49195 0 FreeSerif 160 0 0 0 word693
port 793 nsew
flabel locali -67 -49299 -34 -49266 0 FreeSerif 160 0 0 0 word694
port 794 nsew
flabel locali -67 -49370 -34 -49337 0 FreeSerif 160 0 0 0 word695
port 795 nsew
flabel locali -67 -49441 -34 -49408 0 FreeSerif 160 0 0 0 word696
port 796 nsew
flabel locali -67 -49512 -34 -49479 0 FreeSerif 160 0 0 0 word697
port 797 nsew
flabel locali -67 -49583 -34 -49550 0 FreeSerif 160 0 0 0 word698
port 798 nsew
flabel locali -67 -49654 -34 -49621 0 FreeSerif 160 0 0 0 word699
port 799 nsew
flabel locali -67 -49725 -34 -49692 0 FreeSerif 160 0 0 0 word700
port 800 nsew
flabel locali -67 -49796 -34 -49763 0 FreeSerif 160 0 0 0 word701
port 801 nsew
flabel locali -67 -49867 -34 -49834 0 FreeSerif 160 0 0 0 word702
port 802 nsew
flabel locali -67 -49938 -34 -49905 0 FreeSerif 160 0 0 0 word703
port 803 nsew
flabel locali -67 -50009 -34 -49976 0 FreeSerif 160 0 0 0 word704
port 804 nsew
flabel locali -67 -50080 -34 -50047 0 FreeSerif 160 0 0 0 word705
port 805 nsew
flabel locali -67 -50151 -34 -50118 0 FreeSerif 160 0 0 0 word706
port 806 nsew
flabel locali -67 -50222 -34 -50189 0 FreeSerif 160 0 0 0 word707
port 807 nsew
flabel locali -67 -50293 -34 -50260 0 FreeSerif 160 0 0 0 word708
port 808 nsew
flabel locali -67 -50364 -34 -50331 0 FreeSerif 160 0 0 0 word709
port 809 nsew
flabel locali -67 -50435 -34 -50402 0 FreeSerif 160 0 0 0 word710
port 810 nsew
flabel locali -67 -50506 -34 -50473 0 FreeSerif 160 0 0 0 word711
port 811 nsew
flabel locali -67 -50577 -34 -50544 0 FreeSerif 160 0 0 0 word712
port 812 nsew
flabel locali -67 -50648 -34 -50615 0 FreeSerif 160 0 0 0 word713
port 813 nsew
flabel locali -67 -50719 -34 -50686 0 FreeSerif 160 0 0 0 word714
port 814 nsew
flabel locali -67 -50790 -34 -50757 0 FreeSerif 160 0 0 0 word715
port 815 nsew
flabel locali -67 -50861 -34 -50828 0 FreeSerif 160 0 0 0 word716
port 816 nsew
flabel locali -67 -50932 -34 -50899 0 FreeSerif 160 0 0 0 word717
port 817 nsew
flabel locali -67 -51003 -34 -50970 0 FreeSerif 160 0 0 0 word718
port 818 nsew
flabel locali -67 -51074 -34 -51041 0 FreeSerif 160 0 0 0 word719
port 819 nsew
flabel locali -67 -51145 -34 -51112 0 FreeSerif 160 0 0 0 word720
port 820 nsew
flabel locali -67 -51216 -34 -51183 0 FreeSerif 160 0 0 0 word721
port 821 nsew
flabel locali -67 -51287 -34 -51254 0 FreeSerif 160 0 0 0 word722
port 822 nsew
flabel locali -67 -51358 -34 -51325 0 FreeSerif 160 0 0 0 word723
port 823 nsew
flabel locali -67 -51429 -34 -51396 0 FreeSerif 160 0 0 0 word724
port 824 nsew
flabel locali -67 -51500 -34 -51467 0 FreeSerif 160 0 0 0 word725
port 825 nsew
flabel locali -67 -51571 -34 -51538 0 FreeSerif 160 0 0 0 word726
port 826 nsew
flabel locali -67 -51642 -34 -51609 0 FreeSerif 160 0 0 0 word727
port 827 nsew
flabel locali -67 -51713 -34 -51680 0 FreeSerif 160 0 0 0 word728
port 828 nsew
flabel locali -67 -51784 -34 -51751 0 FreeSerif 160 0 0 0 word729
port 829 nsew
flabel locali -67 -51855 -34 -51822 0 FreeSerif 160 0 0 0 word730
port 830 nsew
flabel locali -67 -51926 -34 -51893 0 FreeSerif 160 0 0 0 word731
port 831 nsew
flabel locali -67 -51997 -34 -51964 0 FreeSerif 160 0 0 0 word732
port 832 nsew
flabel locali -67 -52068 -34 -52035 0 FreeSerif 160 0 0 0 word733
port 833 nsew
flabel locali -67 -52139 -34 -52106 0 FreeSerif 160 0 0 0 word734
port 834 nsew
flabel locali -67 -52210 -34 -52177 0 FreeSerif 160 0 0 0 word735
port 835 nsew
flabel locali -67 -52281 -34 -52248 0 FreeSerif 160 0 0 0 word736
port 836 nsew
flabel locali -67 -52352 -34 -52319 0 FreeSerif 160 0 0 0 word737
port 837 nsew
flabel locali -67 -52423 -34 -52390 0 FreeSerif 160 0 0 0 word738
port 838 nsew
flabel locali -67 -52494 -34 -52461 0 FreeSerif 160 0 0 0 word739
port 839 nsew
flabel locali -67 -52565 -34 -52532 0 FreeSerif 160 0 0 0 word740
port 840 nsew
flabel locali -67 -52636 -34 -52603 0 FreeSerif 160 0 0 0 word741
port 841 nsew
flabel locali -67 -52707 -34 -52674 0 FreeSerif 160 0 0 0 word742
port 842 nsew
flabel locali -67 -52778 -34 -52745 0 FreeSerif 160 0 0 0 word743
port 843 nsew
flabel locali -67 -52849 -34 -52816 0 FreeSerif 160 0 0 0 word744
port 844 nsew
flabel locali -67 -52920 -34 -52887 0 FreeSerif 160 0 0 0 word745
port 845 nsew
flabel locali -67 -52991 -34 -52958 0 FreeSerif 160 0 0 0 word746
port 846 nsew
flabel locali -67 -53062 -34 -53029 0 FreeSerif 160 0 0 0 word747
port 847 nsew
flabel locali -67 -53133 -34 -53100 0 FreeSerif 160 0 0 0 word748
port 848 nsew
flabel locali -67 -53204 -34 -53171 0 FreeSerif 160 0 0 0 word749
port 849 nsew
flabel locali -67 -53275 -34 -53242 0 FreeSerif 160 0 0 0 word750
port 850 nsew
flabel locali -67 -53346 -34 -53313 0 FreeSerif 160 0 0 0 word751
port 851 nsew
flabel locali -67 -53417 -34 -53384 0 FreeSerif 160 0 0 0 word752
port 852 nsew
flabel locali -67 -53488 -34 -53455 0 FreeSerif 160 0 0 0 word753
port 853 nsew
flabel locali -67 -53559 -34 -53526 0 FreeSerif 160 0 0 0 word754
port 854 nsew
flabel locali -67 -53630 -34 -53597 0 FreeSerif 160 0 0 0 word755
port 855 nsew
flabel locali -67 -53701 -34 -53668 0 FreeSerif 160 0 0 0 word756
port 856 nsew
flabel locali -67 -53772 -34 -53739 0 FreeSerif 160 0 0 0 word757
port 857 nsew
flabel locali -67 -53843 -34 -53810 0 FreeSerif 160 0 0 0 word758
port 858 nsew
flabel locali -67 -53914 -34 -53881 0 FreeSerif 160 0 0 0 word759
port 859 nsew
flabel locali -67 -53985 -34 -53952 0 FreeSerif 160 0 0 0 word760
port 860 nsew
flabel locali -67 -54056 -34 -54023 0 FreeSerif 160 0 0 0 word761
port 861 nsew
flabel locali -67 -54127 -34 -54094 0 FreeSerif 160 0 0 0 word762
port 862 nsew
flabel locali -67 -54198 -34 -54165 0 FreeSerif 160 0 0 0 word763
port 863 nsew
flabel locali -67 -54269 -34 -54236 0 FreeSerif 160 0 0 0 word764
port 864 nsew
flabel locali -67 -54340 -34 -54307 0 FreeSerif 160 0 0 0 word765
port 865 nsew
flabel locali -67 -54411 -34 -54378 0 FreeSerif 160 0 0 0 word766
port 866 nsew
flabel locali -67 -54482 -34 -54449 0 FreeSerif 160 0 0 0 word767
port 867 nsew
flabel locali -67 -54553 -34 -54520 0 FreeSerif 160 0 0 0 word768
port 868 nsew
flabel locali -67 -54624 -34 -54591 0 FreeSerif 160 0 0 0 word769
port 869 nsew
flabel locali -67 -54695 -34 -54662 0 FreeSerif 160 0 0 0 word770
port 870 nsew
flabel locali -67 -54766 -34 -54733 0 FreeSerif 160 0 0 0 word771
port 871 nsew
flabel locali -67 -54837 -34 -54804 0 FreeSerif 160 0 0 0 word772
port 872 nsew
flabel locali -67 -54908 -34 -54875 0 FreeSerif 160 0 0 0 word773
port 873 nsew
flabel locali -67 -54979 -34 -54946 0 FreeSerif 160 0 0 0 word774
port 874 nsew
flabel locali -67 -55050 -34 -55017 0 FreeSerif 160 0 0 0 word775
port 875 nsew
flabel locali -67 -55121 -34 -55088 0 FreeSerif 160 0 0 0 word776
port 876 nsew
flabel locali -67 -55192 -34 -55159 0 FreeSerif 160 0 0 0 word777
port 877 nsew
flabel locali -67 -55263 -34 -55230 0 FreeSerif 160 0 0 0 word778
port 878 nsew
flabel locali -67 -55334 -34 -55301 0 FreeSerif 160 0 0 0 word779
port 879 nsew
flabel locali -67 -55405 -34 -55372 0 FreeSerif 160 0 0 0 word780
port 880 nsew
flabel locali -67 -55476 -34 -55443 0 FreeSerif 160 0 0 0 word781
port 881 nsew
flabel locali -67 -55547 -34 -55514 0 FreeSerif 160 0 0 0 word782
port 882 nsew
flabel locali -67 -55618 -34 -55585 0 FreeSerif 160 0 0 0 word783
port 883 nsew
flabel locali -67 -55689 -34 -55656 0 FreeSerif 160 0 0 0 word784
port 884 nsew
flabel locali -67 -55760 -34 -55727 0 FreeSerif 160 0 0 0 word785
port 885 nsew
flabel locali -67 -55831 -34 -55798 0 FreeSerif 160 0 0 0 word786
port 886 nsew
flabel locali -67 -55902 -34 -55869 0 FreeSerif 160 0 0 0 word787
port 887 nsew
flabel locali -67 -55973 -34 -55940 0 FreeSerif 160 0 0 0 word788
port 888 nsew
flabel locali -67 -56044 -34 -56011 0 FreeSerif 160 0 0 0 word789
port 889 nsew
flabel locali -67 -56115 -34 -56082 0 FreeSerif 160 0 0 0 word790
port 890 nsew
flabel locali -67 -56186 -34 -56153 0 FreeSerif 160 0 0 0 word791
port 891 nsew
flabel locali -67 -56257 -34 -56224 0 FreeSerif 160 0 0 0 word792
port 892 nsew
flabel locali -67 -56328 -34 -56295 0 FreeSerif 160 0 0 0 word793
port 893 nsew
flabel locali -67 -56399 -34 -56366 0 FreeSerif 160 0 0 0 word794
port 894 nsew
flabel locali -67 -56470 -34 -56437 0 FreeSerif 160 0 0 0 word795
port 895 nsew
flabel locali -67 -56541 -34 -56508 0 FreeSerif 160 0 0 0 word796
port 896 nsew
flabel locali -67 -56612 -34 -56579 0 FreeSerif 160 0 0 0 word797
port 897 nsew
flabel locali -67 -56683 -34 -56650 0 FreeSerif 160 0 0 0 word798
port 898 nsew
flabel locali -67 -56754 -34 -56721 0 FreeSerif 160 0 0 0 word799
port 899 nsew
flabel locali -67 -56825 -34 -56792 0 FreeSerif 160 0 0 0 word800
port 900 nsew
flabel locali -67 -56896 -34 -56863 0 FreeSerif 160 0 0 0 word801
port 901 nsew
flabel locali -67 -56967 -34 -56934 0 FreeSerif 160 0 0 0 word802
port 902 nsew
flabel locali -67 -57038 -34 -57005 0 FreeSerif 160 0 0 0 word803
port 903 nsew
flabel locali -67 -57109 -34 -57076 0 FreeSerif 160 0 0 0 word804
port 904 nsew
flabel locali -67 -57180 -34 -57147 0 FreeSerif 160 0 0 0 word805
port 905 nsew
flabel locali -67 -57251 -34 -57218 0 FreeSerif 160 0 0 0 word806
port 906 nsew
flabel locali -67 -57322 -34 -57289 0 FreeSerif 160 0 0 0 word807
port 907 nsew
flabel locali -67 -57393 -34 -57360 0 FreeSerif 160 0 0 0 word808
port 908 nsew
flabel locali -67 -57464 -34 -57431 0 FreeSerif 160 0 0 0 word809
port 909 nsew
flabel locali -67 -57535 -34 -57502 0 FreeSerif 160 0 0 0 word810
port 910 nsew
flabel locali -67 -57606 -34 -57573 0 FreeSerif 160 0 0 0 word811
port 911 nsew
flabel locali -67 -57677 -34 -57644 0 FreeSerif 160 0 0 0 word812
port 912 nsew
flabel locali -67 -57748 -34 -57715 0 FreeSerif 160 0 0 0 word813
port 913 nsew
flabel locali -67 -57819 -34 -57786 0 FreeSerif 160 0 0 0 word814
port 914 nsew
flabel locali -67 -57890 -34 -57857 0 FreeSerif 160 0 0 0 word815
port 915 nsew
flabel locali -67 -57961 -34 -57928 0 FreeSerif 160 0 0 0 word816
port 916 nsew
flabel locali -67 -58032 -34 -57999 0 FreeSerif 160 0 0 0 word817
port 917 nsew
flabel locali -67 -58103 -34 -58070 0 FreeSerif 160 0 0 0 word818
port 918 nsew
flabel locali -67 -58174 -34 -58141 0 FreeSerif 160 0 0 0 word819
port 919 nsew
flabel locali -67 -58245 -34 -58212 0 FreeSerif 160 0 0 0 word820
port 920 nsew
flabel locali -67 -58316 -34 -58283 0 FreeSerif 160 0 0 0 word821
port 921 nsew
flabel locali -67 -58387 -34 -58354 0 FreeSerif 160 0 0 0 word822
port 922 nsew
flabel locali -67 -58458 -34 -58425 0 FreeSerif 160 0 0 0 word823
port 923 nsew
flabel locali -67 -58529 -34 -58496 0 FreeSerif 160 0 0 0 word824
port 924 nsew
flabel locali -67 -58600 -34 -58567 0 FreeSerif 160 0 0 0 word825
port 925 nsew
flabel locali -67 -58671 -34 -58638 0 FreeSerif 160 0 0 0 word826
port 926 nsew
flabel locali -67 -58742 -34 -58709 0 FreeSerif 160 0 0 0 word827
port 927 nsew
flabel locali -67 -58813 -34 -58780 0 FreeSerif 160 0 0 0 word828
port 928 nsew
flabel locali -67 -58884 -34 -58851 0 FreeSerif 160 0 0 0 word829
port 929 nsew
flabel locali -67 -58955 -34 -58922 0 FreeSerif 160 0 0 0 word830
port 930 nsew
flabel locali -67 -59026 -34 -58993 0 FreeSerif 160 0 0 0 word831
port 931 nsew
flabel locali -67 -59097 -34 -59064 0 FreeSerif 160 0 0 0 word832
port 932 nsew
flabel locali -67 -59168 -34 -59135 0 FreeSerif 160 0 0 0 word833
port 933 nsew
flabel locali -67 -59239 -34 -59206 0 FreeSerif 160 0 0 0 word834
port 934 nsew
flabel locali -67 -59310 -34 -59277 0 FreeSerif 160 0 0 0 word835
port 935 nsew
flabel locali -67 -59381 -34 -59348 0 FreeSerif 160 0 0 0 word836
port 936 nsew
flabel locali -67 -59452 -34 -59419 0 FreeSerif 160 0 0 0 word837
port 937 nsew
flabel locali -67 -59523 -34 -59490 0 FreeSerif 160 0 0 0 word838
port 938 nsew
flabel locali -67 -59594 -34 -59561 0 FreeSerif 160 0 0 0 word839
port 939 nsew
flabel locali -67 -59665 -34 -59632 0 FreeSerif 160 0 0 0 word840
port 940 nsew
flabel locali -67 -59736 -34 -59703 0 FreeSerif 160 0 0 0 word841
port 941 nsew
flabel locali -67 -59807 -34 -59774 0 FreeSerif 160 0 0 0 word842
port 942 nsew
flabel locali -67 -59878 -34 -59845 0 FreeSerif 160 0 0 0 word843
port 943 nsew
flabel locali -67 -59949 -34 -59916 0 FreeSerif 160 0 0 0 word844
port 944 nsew
flabel locali -67 -60020 -34 -59987 0 FreeSerif 160 0 0 0 word845
port 945 nsew
flabel locali -67 -60091 -34 -60058 0 FreeSerif 160 0 0 0 word846
port 946 nsew
flabel locali -67 -60162 -34 -60129 0 FreeSerif 160 0 0 0 word847
port 947 nsew
flabel locali -67 -60233 -34 -60200 0 FreeSerif 160 0 0 0 word848
port 948 nsew
flabel locali -67 -60304 -34 -60271 0 FreeSerif 160 0 0 0 word849
port 949 nsew
flabel locali -67 -60375 -34 -60342 0 FreeSerif 160 0 0 0 word850
port 950 nsew
flabel locali -67 -60446 -34 -60413 0 FreeSerif 160 0 0 0 word851
port 951 nsew
flabel locali -67 -60517 -34 -60484 0 FreeSerif 160 0 0 0 word852
port 952 nsew
flabel locali -67 -60588 -34 -60555 0 FreeSerif 160 0 0 0 word853
port 953 nsew
flabel locali -67 -60659 -34 -60626 0 FreeSerif 160 0 0 0 word854
port 954 nsew
flabel locali -67 -60730 -34 -60697 0 FreeSerif 160 0 0 0 word855
port 955 nsew
flabel locali -67 -60801 -34 -60768 0 FreeSerif 160 0 0 0 word856
port 956 nsew
flabel locali -67 -60872 -34 -60839 0 FreeSerif 160 0 0 0 word857
port 957 nsew
flabel locali -67 -60943 -34 -60910 0 FreeSerif 160 0 0 0 word858
port 958 nsew
flabel locali -67 -61014 -34 -60981 0 FreeSerif 160 0 0 0 word859
port 959 nsew
flabel locali -67 -61085 -34 -61052 0 FreeSerif 160 0 0 0 word860
port 960 nsew
flabel locali -67 -61156 -34 -61123 0 FreeSerif 160 0 0 0 word861
port 961 nsew
flabel locali -67 -61227 -34 -61194 0 FreeSerif 160 0 0 0 word862
port 962 nsew
flabel locali -67 -61298 -34 -61265 0 FreeSerif 160 0 0 0 word863
port 963 nsew
flabel locali -67 -61369 -34 -61336 0 FreeSerif 160 0 0 0 word864
port 964 nsew
flabel locali -67 -61440 -34 -61407 0 FreeSerif 160 0 0 0 word865
port 965 nsew
flabel locali -67 -61511 -34 -61478 0 FreeSerif 160 0 0 0 word866
port 966 nsew
flabel locali -67 -61582 -34 -61549 0 FreeSerif 160 0 0 0 word867
port 967 nsew
flabel locali -67 -61653 -34 -61620 0 FreeSerif 160 0 0 0 word868
port 968 nsew
flabel locali -67 -61724 -34 -61691 0 FreeSerif 160 0 0 0 word869
port 969 nsew
flabel locali -67 -61795 -34 -61762 0 FreeSerif 160 0 0 0 word870
port 970 nsew
flabel locali -67 -61866 -34 -61833 0 FreeSerif 160 0 0 0 word871
port 971 nsew
flabel locali -67 -61937 -34 -61904 0 FreeSerif 160 0 0 0 word872
port 972 nsew
flabel locali -67 -62008 -34 -61975 0 FreeSerif 160 0 0 0 word873
port 973 nsew
flabel locali -67 -62079 -34 -62046 0 FreeSerif 160 0 0 0 word874
port 974 nsew
flabel locali -67 -62150 -34 -62117 0 FreeSerif 160 0 0 0 word875
port 975 nsew
flabel locali -67 -62221 -34 -62188 0 FreeSerif 160 0 0 0 word876
port 976 nsew
flabel locali -67 -62292 -34 -62259 0 FreeSerif 160 0 0 0 word877
port 977 nsew
flabel locali -67 -62363 -34 -62330 0 FreeSerif 160 0 0 0 word878
port 978 nsew
flabel locali -67 -62434 -34 -62401 0 FreeSerif 160 0 0 0 word879
port 979 nsew
flabel locali -67 -62505 -34 -62472 0 FreeSerif 160 0 0 0 word880
port 980 nsew
flabel locali -67 -62576 -34 -62543 0 FreeSerif 160 0 0 0 word881
port 981 nsew
flabel locali -67 -62647 -34 -62614 0 FreeSerif 160 0 0 0 word882
port 982 nsew
flabel locali -67 -62718 -34 -62685 0 FreeSerif 160 0 0 0 word883
port 983 nsew
flabel locali -67 -62789 -34 -62756 0 FreeSerif 160 0 0 0 word884
port 984 nsew
flabel locali -67 -62860 -34 -62827 0 FreeSerif 160 0 0 0 word885
port 985 nsew
flabel locali -67 -62931 -34 -62898 0 FreeSerif 160 0 0 0 word886
port 986 nsew
flabel locali -67 -63002 -34 -62969 0 FreeSerif 160 0 0 0 word887
port 987 nsew
flabel locali -67 -63073 -34 -63040 0 FreeSerif 160 0 0 0 word888
port 988 nsew
flabel locali -67 -63144 -34 -63111 0 FreeSerif 160 0 0 0 word889
port 989 nsew
flabel locali -67 -63215 -34 -63182 0 FreeSerif 160 0 0 0 word890
port 990 nsew
flabel locali -67 -63286 -34 -63253 0 FreeSerif 160 0 0 0 word891
port 991 nsew
flabel locali -67 -63357 -34 -63324 0 FreeSerif 160 0 0 0 word892
port 992 nsew
flabel locali -67 -63428 -34 -63395 0 FreeSerif 160 0 0 0 word893
port 993 nsew
flabel locali -67 -63499 -34 -63466 0 FreeSerif 160 0 0 0 word894
port 994 nsew
flabel locali -67 -63570 -34 -63537 0 FreeSerif 160 0 0 0 word895
port 995 nsew
flabel locali -67 -63641 -34 -63608 0 FreeSerif 160 0 0 0 word896
port 996 nsew
flabel locali -67 -63712 -34 -63679 0 FreeSerif 160 0 0 0 word897
port 997 nsew
flabel locali -67 -63783 -34 -63750 0 FreeSerif 160 0 0 0 word898
port 998 nsew
flabel locali -67 -63854 -34 -63821 0 FreeSerif 160 0 0 0 word899
port 999 nsew
flabel locali -67 -63925 -34 -63892 0 FreeSerif 160 0 0 0 word900
port 1000 nsew
flabel locali -67 -63996 -34 -63963 0 FreeSerif 160 0 0 0 word901
port 1001 nsew
flabel locali -67 -64067 -34 -64034 0 FreeSerif 160 0 0 0 word902
port 1002 nsew
flabel locali -67 -64138 -34 -64105 0 FreeSerif 160 0 0 0 word903
port 1003 nsew
flabel locali -67 -64209 -34 -64176 0 FreeSerif 160 0 0 0 word904
port 1004 nsew
flabel locali -67 -64280 -34 -64247 0 FreeSerif 160 0 0 0 word905
port 1005 nsew
flabel locali -67 -64351 -34 -64318 0 FreeSerif 160 0 0 0 word906
port 1006 nsew
flabel locali -67 -64422 -34 -64389 0 FreeSerif 160 0 0 0 word907
port 1007 nsew
flabel locali -67 -64493 -34 -64460 0 FreeSerif 160 0 0 0 word908
port 1008 nsew
flabel locali -67 -64564 -34 -64531 0 FreeSerif 160 0 0 0 word909
port 1009 nsew
flabel locali -67 -64635 -34 -64602 0 FreeSerif 160 0 0 0 word910
port 1010 nsew
flabel locali -67 -64706 -34 -64673 0 FreeSerif 160 0 0 0 word911
port 1011 nsew
flabel locali -67 -64777 -34 -64744 0 FreeSerif 160 0 0 0 word912
port 1012 nsew
flabel locali -67 -64848 -34 -64815 0 FreeSerif 160 0 0 0 word913
port 1013 nsew
flabel locali -67 -64919 -34 -64886 0 FreeSerif 160 0 0 0 word914
port 1014 nsew
flabel locali -67 -64990 -34 -64957 0 FreeSerif 160 0 0 0 word915
port 1015 nsew
flabel locali -67 -65061 -34 -65028 0 FreeSerif 160 0 0 0 word916
port 1016 nsew
flabel locali -67 -65132 -34 -65099 0 FreeSerif 160 0 0 0 word917
port 1017 nsew
flabel locali -67 -65203 -34 -65170 0 FreeSerif 160 0 0 0 word918
port 1018 nsew
flabel locali -67 -65274 -34 -65241 0 FreeSerif 160 0 0 0 word919
port 1019 nsew
flabel locali -67 -65345 -34 -65312 0 FreeSerif 160 0 0 0 word920
port 1020 nsew
flabel locali -67 -65416 -34 -65383 0 FreeSerif 160 0 0 0 word921
port 1021 nsew
flabel locali -67 -65487 -34 -65454 0 FreeSerif 160 0 0 0 word922
port 1022 nsew
flabel locali -67 -65558 -34 -65525 0 FreeSerif 160 0 0 0 word923
port 1023 nsew
flabel locali -67 -65629 -34 -65596 0 FreeSerif 160 0 0 0 word924
port 1024 nsew
flabel locali -67 -65700 -34 -65667 0 FreeSerif 160 0 0 0 word925
port 1025 nsew
flabel locali -67 -65771 -34 -65738 0 FreeSerif 160 0 0 0 word926
port 1026 nsew
flabel locali -67 -65842 -34 -65809 0 FreeSerif 160 0 0 0 word927
port 1027 nsew
flabel locali -67 -65913 -34 -65880 0 FreeSerif 160 0 0 0 word928
port 1028 nsew
flabel locali -67 -65984 -34 -65951 0 FreeSerif 160 0 0 0 word929
port 1029 nsew
flabel locali -67 -66055 -34 -66022 0 FreeSerif 160 0 0 0 word930
port 1030 nsew
flabel locali -67 -66126 -34 -66093 0 FreeSerif 160 0 0 0 word931
port 1031 nsew
flabel locali -67 -66197 -34 -66164 0 FreeSerif 160 0 0 0 word932
port 1032 nsew
flabel locali -67 -66268 -34 -66235 0 FreeSerif 160 0 0 0 word933
port 1033 nsew
flabel locali -67 -66339 -34 -66306 0 FreeSerif 160 0 0 0 word934
port 1034 nsew
flabel locali -67 -66410 -34 -66377 0 FreeSerif 160 0 0 0 word935
port 1035 nsew
flabel locali -67 -66481 -34 -66448 0 FreeSerif 160 0 0 0 word936
port 1036 nsew
flabel locali -67 -66552 -34 -66519 0 FreeSerif 160 0 0 0 word937
port 1037 nsew
flabel locali -67 -66623 -34 -66590 0 FreeSerif 160 0 0 0 word938
port 1038 nsew
flabel locali -67 -66694 -34 -66661 0 FreeSerif 160 0 0 0 word939
port 1039 nsew
flabel locali -67 -66765 -34 -66732 0 FreeSerif 160 0 0 0 word940
port 1040 nsew
flabel locali -67 -66836 -34 -66803 0 FreeSerif 160 0 0 0 word941
port 1041 nsew
flabel locali -67 -66907 -34 -66874 0 FreeSerif 160 0 0 0 word942
port 1042 nsew
flabel locali -67 -66978 -34 -66945 0 FreeSerif 160 0 0 0 word943
port 1043 nsew
flabel locali -67 -67049 -34 -67016 0 FreeSerif 160 0 0 0 word944
port 1044 nsew
flabel locali -67 -67120 -34 -67087 0 FreeSerif 160 0 0 0 word945
port 1045 nsew
flabel locali -67 -67191 -34 -67158 0 FreeSerif 160 0 0 0 word946
port 1046 nsew
flabel locali -67 -67262 -34 -67229 0 FreeSerif 160 0 0 0 word947
port 1047 nsew
flabel locali -67 -67333 -34 -67300 0 FreeSerif 160 0 0 0 word948
port 1048 nsew
flabel locali -67 -67404 -34 -67371 0 FreeSerif 160 0 0 0 word949
port 1049 nsew
flabel locali -67 -67475 -34 -67442 0 FreeSerif 160 0 0 0 word950
port 1050 nsew
flabel locali -67 -67546 -34 -67513 0 FreeSerif 160 0 0 0 word951
port 1051 nsew
flabel locali -67 -67617 -34 -67584 0 FreeSerif 160 0 0 0 word952
port 1052 nsew
flabel locali -67 -67688 -34 -67655 0 FreeSerif 160 0 0 0 word953
port 1053 nsew
flabel locali -67 -67759 -34 -67726 0 FreeSerif 160 0 0 0 word954
port 1054 nsew
flabel locali -67 -67830 -34 -67797 0 FreeSerif 160 0 0 0 word955
port 1055 nsew
flabel locali -67 -67901 -34 -67868 0 FreeSerif 160 0 0 0 word956
port 1056 nsew
flabel locali -67 -67972 -34 -67939 0 FreeSerif 160 0 0 0 word957
port 1057 nsew
flabel locali -67 -68043 -34 -68010 0 FreeSerif 160 0 0 0 word958
port 1058 nsew
flabel locali -67 -68114 -34 -68081 0 FreeSerif 160 0 0 0 word959
port 1059 nsew
flabel locali -67 -68185 -34 -68152 0 FreeSerif 160 0 0 0 word960
port 1060 nsew
flabel locali -67 -68256 -34 -68223 0 FreeSerif 160 0 0 0 word961
port 1061 nsew
flabel locali -67 -68327 -34 -68294 0 FreeSerif 160 0 0 0 word962
port 1062 nsew
flabel locali -67 -68398 -34 -68365 0 FreeSerif 160 0 0 0 word963
port 1063 nsew
flabel locali -67 -68469 -34 -68436 0 FreeSerif 160 0 0 0 word964
port 1064 nsew
flabel locali -67 -68540 -34 -68507 0 FreeSerif 160 0 0 0 word965
port 1065 nsew
flabel locali -67 -68611 -34 -68578 0 FreeSerif 160 0 0 0 word966
port 1066 nsew
flabel locali -67 -68682 -34 -68649 0 FreeSerif 160 0 0 0 word967
port 1067 nsew
flabel locali -67 -68753 -34 -68720 0 FreeSerif 160 0 0 0 word968
port 1068 nsew
flabel locali -67 -68824 -34 -68791 0 FreeSerif 160 0 0 0 word969
port 1069 nsew
flabel locali -67 -68895 -34 -68862 0 FreeSerif 160 0 0 0 word970
port 1070 nsew
flabel locali -67 -68966 -34 -68933 0 FreeSerif 160 0 0 0 word971
port 1071 nsew
flabel locali -67 -69037 -34 -69004 0 FreeSerif 160 0 0 0 word972
port 1072 nsew
flabel locali -67 -69108 -34 -69075 0 FreeSerif 160 0 0 0 word973
port 1073 nsew
flabel locali -67 -69179 -34 -69146 0 FreeSerif 160 0 0 0 word974
port 1074 nsew
flabel locali -67 -69250 -34 -69217 0 FreeSerif 160 0 0 0 word975
port 1075 nsew
flabel locali -67 -69321 -34 -69288 0 FreeSerif 160 0 0 0 word976
port 1076 nsew
flabel locali -67 -69392 -34 -69359 0 FreeSerif 160 0 0 0 word977
port 1077 nsew
flabel locali -67 -69463 -34 -69430 0 FreeSerif 160 0 0 0 word978
port 1078 nsew
flabel locali -67 -69534 -34 -69501 0 FreeSerif 160 0 0 0 word979
port 1079 nsew
flabel locali -67 -69605 -34 -69572 0 FreeSerif 160 0 0 0 word980
port 1080 nsew
flabel locali -67 -69676 -34 -69643 0 FreeSerif 160 0 0 0 word981
port 1081 nsew
flabel locali -67 -69747 -34 -69714 0 FreeSerif 160 0 0 0 word982
port 1082 nsew
flabel locali -67 -69818 -34 -69785 0 FreeSerif 160 0 0 0 word983
port 1083 nsew
flabel locali -67 -69889 -34 -69856 0 FreeSerif 160 0 0 0 word984
port 1084 nsew
flabel locali -67 -69960 -34 -69927 0 FreeSerif 160 0 0 0 word985
port 1085 nsew
flabel locali -67 -70031 -34 -69998 0 FreeSerif 160 0 0 0 word986
port 1086 nsew
flabel locali -67 -70102 -34 -70069 0 FreeSerif 160 0 0 0 word987
port 1087 nsew
flabel locali -67 -70173 -34 -70140 0 FreeSerif 160 0 0 0 word988
port 1088 nsew
flabel locali -67 -70244 -34 -70211 0 FreeSerif 160 0 0 0 word989
port 1089 nsew
flabel locali -67 -70315 -34 -70282 0 FreeSerif 160 0 0 0 word990
port 1090 nsew
flabel locali -67 -70386 -34 -70353 0 FreeSerif 160 0 0 0 word991
port 1091 nsew
flabel locali -67 -70457 -34 -70424 0 FreeSerif 160 0 0 0 word992
port 1092 nsew
flabel locali -67 -70528 -34 -70495 0 FreeSerif 160 0 0 0 word993
port 1093 nsew
flabel locali -67 -70599 -34 -70566 0 FreeSerif 160 0 0 0 word994
port 1094 nsew
flabel locali -67 -70670 -34 -70637 0 FreeSerif 160 0 0 0 word995
port 1095 nsew
flabel locali -67 -70741 -34 -70708 0 FreeSerif 160 0 0 0 word996
port 1096 nsew
flabel locali -67 -70812 -34 -70779 0 FreeSerif 160 0 0 0 word997
port 1097 nsew
flabel locali -67 -70883 -34 -70850 0 FreeSerif 160 0 0 0 word998
port 1098 nsew
flabel locali -67 -70954 -34 -70921 0 FreeSerif 160 0 0 0 word999
port 1099 nsew
flabel locali -67 -71025 -34 -70992 0 FreeSerif 160 0 0 0 word1000
port 1100 nsew
flabel locali -67 -71096 -34 -71063 0 FreeSerif 160 0 0 0 word1001
port 1101 nsew
flabel locali -67 -71167 -34 -71134 0 FreeSerif 160 0 0 0 word1002
port 1102 nsew
flabel locali -67 -71238 -34 -71205 0 FreeSerif 160 0 0 0 word1003
port 1103 nsew
flabel locali -67 -71309 -34 -71276 0 FreeSerif 160 0 0 0 word1004
port 1104 nsew
flabel locali -67 -71380 -34 -71347 0 FreeSerif 160 0 0 0 word1005
port 1105 nsew
flabel locali -67 -71451 -34 -71418 0 FreeSerif 160 0 0 0 word1006
port 1106 nsew
flabel locali -67 -71522 -34 -71489 0 FreeSerif 160 0 0 0 word1007
port 1107 nsew
flabel locali -67 -71593 -34 -71560 0 FreeSerif 160 0 0 0 word1008
port 1108 nsew
flabel locali -67 -71664 -34 -71631 0 FreeSerif 160 0 0 0 word1009
port 1109 nsew
flabel locali -67 -71735 -34 -71702 0 FreeSerif 160 0 0 0 word1010
port 1110 nsew
flabel locali -67 -71806 -34 -71773 0 FreeSerif 160 0 0 0 word1011
port 1111 nsew
flabel locali -67 -71877 -34 -71844 0 FreeSerif 160 0 0 0 word1012
port 1112 nsew
flabel locali -67 -71948 -34 -71915 0 FreeSerif 160 0 0 0 word1013
port 1113 nsew
flabel locali -67 -72019 -34 -71986 0 FreeSerif 160 0 0 0 word1014
port 1114 nsew
flabel locali -67 -72090 -34 -72057 0 FreeSerif 160 0 0 0 word1015
port 1115 nsew
flabel locali -67 -72161 -34 -72128 0 FreeSerif 160 0 0 0 word1016
port 1116 nsew
flabel locali -67 -72232 -34 -72199 0 FreeSerif 160 0 0 0 word1017
port 1117 nsew
flabel locali -67 -72303 -34 -72270 0 FreeSerif 160 0 0 0 word1018
port 1118 nsew
flabel locali -67 -72374 -34 -72341 0 FreeSerif 160 0 0 0 word1019
port 1119 nsew
flabel locali -67 -72445 -34 -72412 0 FreeSerif 160 0 0 0 word1020
port 1120 nsew
flabel locali -67 -72516 -34 -72483 0 FreeSerif 160 0 0 0 word1021
port 1121 nsew
flabel locali -67 -72587 -34 -72554 0 FreeSerif 160 0 0 0 word1022
port 1122 nsew
flabel locali -67 -72658 -34 -72625 0 FreeSerif 160 0 0 0 word1023
port 1123 nsew
flabel locali 0 -72737 33 -72704 0 FreeSerif 160 0 0 0 Y7
port 1124 nsew
flabel locali 166 -72737 199 -72704 0 FreeSerif 160 0 0 0 Y6
port 1125 nsew
flabel locali 249 -72737 282 -72704 0 FreeSerif 160 0 0 0 Y5
port 1126 nsew
flabel locali 415 -72737 448 -72704 0 FreeSerif 160 0 0 0 Y4
port 1127 nsew
flabel locali 498 -72737 531 -72704 0 FreeSerif 160 0 0 0 Y3
port 1128 nsew
flabel locali 664 -72737 697 -72704 0 FreeSerif 160 0 0 0 Y2
port 1129 nsew
flabel locali 747 -72737 780 -72704 0 FreeSerif 160 0 0 0 Y1
port 1130 nsew
flabel locali 913 -72737 946 -72704 0 FreeSerif 160 0 0 0 Y0
port 1131 nsew
flabel locali -27 69 973 117 0 FreeSerif 160 0 0 0 GND!
port 1132 nsew
flabel locali -25 244 971 292 0 FreeSerif 160 0 0 0 VDD!
port 1133 nsew
<< end >>