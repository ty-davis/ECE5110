* NGSPICE file created from memory_out.ext - technology: sky130A

*.subckt memory_out word0 word1 word2 word3 word4 word5 word6 word7 word8 word9 word10
+ word11 word12 word13 word14 word15 word16 word17 word18 word19 word20 word21 word22
+ word23 word24 word25 word26 word27 word28 word29 word30 word31 word32 word33 word34
+ word35 word36 word37 word38 word39 word40 word41 word42 word43 word44 word45 word46
+ word47 word48 word49 word50 word51 word52 word53 word54 word55 word56 word57 word58
+ word59 word60 word61 word62 word63 word64 word65 word66 word67 word68 word69 word70
+ word71 word72 word73 word74 word75 word76 word77 word78 word79 word80 word81 word82
+ word83 word84 word85 word86 word87 word88 word89 word90 word91 word92 word93 word94
+ word95 word96 word97 word98 word99 word100 word101 word102 word103 word104 word105
+ word106 word107 word108 word109 word110 word111 word112 word113 word114 word115
+ word116 word117 word118 word119 word120 word121 word122 word123 word124 word125
+ word126 word127 Y7 Y6 Y5 Y4 Y3 Y2 Y1 Y0 GND VDD
X0 GND word73 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1 Y7 word52 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2 GND word49 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3 GND word107 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X4 Y2 word66 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X5 Y4 word46 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X6 Y5 word106 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X7 GND word99 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X8 Y2 word48 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X9 GND word33 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X10 GND word35 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X11 GND word17 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X12 Y6 word102 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X13 Y1 word30 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X14 GND word115 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X15 GND word93 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X16 VDD GND Y5 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X17 GND word43 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X18 GND word71 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X19 Y0 word24 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X20 Y2 word110 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X21 Y0 word70 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X22 GND word59 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X23 GND word57 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X24 GND word39 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X25 GND word41 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X26 Y3 word126 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X27 GND word93 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X28 GND word99 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X29 GND word21 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X30 GND word19 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X31 Y1 word112 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X32 Y4 word48 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X33 Y1 word92 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X34 GND word61 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X35 Y1 word50 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X36 Y3 word30 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X37 Y0 word110 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X38 Y4 word106 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X39 Y7 word42 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X40 GND word115 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X41 GND word121 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X42 Y0 word26 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X43 Y2 word112 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X44 GND word103 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X45 GND word59 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X46 Y6 word58 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X47 Y2 word56 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X48 GND word41 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X49 GND word25 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X50 Y5 word28 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X51 Y2 word92 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X52 Y6 word110 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X53 GND word71 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X54 GND word23 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X55 Y3 word108 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X56 GND word101 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X57 Y6 word20 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X58 GND word19 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X59 GND word79 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X60 GND word51 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X61 GND word35 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X62 GND word121 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X63 GND word17 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X64 Y7 word106 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X65 GND word103 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X66 GND word65 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X67 GND word63 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X68 Y1 word52 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X69 Y3 word50 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X70 GND word49 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X71 Y0 word112 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X72 Y7 word16 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X73 Y4 word108 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X74 Y1 word74 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X75 GND word29 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X76 Y0 word92 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X77 GND word117 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X78 Y4 word56 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X79 GND word27 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X80 GND word43 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X81 Y6 word112 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X82 GND word23 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X83 GND word121 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X84 Y6 word40 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X85 GND word103 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X86 Y6 word92 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X87 GND word53 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X88 Y2 word74 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X89 Y0 word34 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X90 GND word21 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X91 Y7 word108 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X92 Y3 word90 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X93 GND word69 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X94 GND word67 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X95 Y3 word52 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X96 GND word49 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X97 Y5 word36 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X98 GND word121 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X99 Y5 word18 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X100 GND word79 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X101 GND word125 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X102 GND word103 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X103 VDD GND Y7 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X104 Y1 word76 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X105 GND word31 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X106 Y5 word72 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X107 GND word25 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X108 Y0 word28 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X109 Y5 word118 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X110 GND word47 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X111 GND word111 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X112 Y1 word60 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X113 Y2 word58 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X114 GND word43 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X115 Y1 word42 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X116 Y0 word74 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X117 Y7 word24 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X118 GND word85 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X119 Y0 word54 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X120 Y2 word76 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X121 GND word21 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X122 Y6 word22 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X123 Y2 word20 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X124 GND word67 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X125 Y6 word74 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X126 GND word51 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X127 Y3 word72 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X128 GND word111 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X129 Y7 word90 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X130 VDD GND Y2 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X131 GND word85 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X132 VDD GND Y3 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X133 GND word45 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X134 Y1 word122 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X135 GND word27 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X136 GND word29 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X137 Y1 word16 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X138 Y1 word62 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X139 Y3 word60 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X140 Y4 word58 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X141 Y3 word42 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X142 Y5 word44 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X143 Y0 word76 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X144 Y7 word26 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X145 GND word111 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X146 Y4 word72 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X147 Y4 word118 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X148 Y1 word84 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X149 GND word39 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X150 GND word81 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X151 Y2 word40 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X152 Y4 word20 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X153 Y5 word80 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X154 Y0 word36 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X155 Y2 word122 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X156 Y0 word18 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X157 Y6 word76 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X158 GND word85 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X159 GND word51 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X160 GND word83 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X161 GND word53 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X162 GND word109 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X163 GND word17 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X164 Y1 word78 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X165 GND word47 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X166 Y2 word84 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X167 GND word75 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X168 GND word29 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X169 Y6 word30 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X170 GND word31 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X171 Y7 word118 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X172 Y3 word16 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X173 Y3 word62 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X174 GND word113 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X175 Y3 word80 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X176 Y0 word122 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X177 GND word59 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X178 GND word83 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X179 Y4 word40 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X180 Y5 word100 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X181 Y0 word38 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X182 Y2 word78 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X183 GND word75 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X184 Y2 word22 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X185 Y1 word24 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X186 GND word109 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X187 Y1 word70 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X188 Y2 word68 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X189 Y0 word84 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X190 GND word53 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X191 Y6 word122 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X192 Y4 word80 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X193 GND word113 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X194 GND word95 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X195 GND word89 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X196 GND word77 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X197 Y6 word50 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X198 GND word31 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X199 GND word33 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X200 Y0 word44 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X201 Y5 word48 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X202 GND word91 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X203 Y3 word82 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X204 GND word61 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X205 Y0 word78 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X206 GND word75 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X207 Y7 word28 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X208 GND word113 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X209 GND word25 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X210 GND word95 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X211 Y1 word86 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X212 GND word55 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X213 GND word39 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X214 GND word77 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X215 Y4 word22 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X216 GND word23 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X217 Y3 word24 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X218 Y1 word26 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X219 Y3 word70 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X220 Y4 word68 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X221 GND word57 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X222 Y6 word78 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X223 GND word75 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X224 Y7 word54 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X225 GND word109 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X226 GND word97 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X227 GND word91 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X228 GND word49 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X229 GND word93 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X230 GND word19 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X231 Y2 word86 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X232 GND word35 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X233 Y0 word46 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X234 Y2 word30 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X235 GND word17 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X236 Y3 word102 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X237 GND word95 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X238 GND word63 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X239 GND word61 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X240 GND word77 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X241 GND word45 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X242 GND word27 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X243 Y1 word88 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X244 GND word59 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X245 Y7 word82 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X246 GND word41 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X247 Y3 word26 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X248 GND word37 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X249 GND word95 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X250 Y5 word56 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X251 GND word77 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X252 Y0 word86 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X253 VDD GND Y0 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X254 Y5 word110 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X255 Y7 word18 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X256 Y1 word94 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X257 Y0 word66 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X258 Y2 word88 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X259 Y2 word50 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X260 Y0 word48 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X261 Y4 word30 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X262 Y1 word34 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X263 GND word35 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X264 GND word17 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X265 GND word119 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X266 GND word63 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X267 GND word47 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X268 GND word123 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X269 GND word101 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X270 Y2 word94 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X271 GND word57 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X272 GND word23 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X273 GND word25 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X274 Y1 word28 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X275 GND word119 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X276 Y0 word88 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X277 GND word99 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X278 GND word19 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X279 Y5 word112 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X280 VDD GND Y1 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X281 GND word93 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X282 Y1 word54 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X283 Y2 word52 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X284 GND word51 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X285 Y4 word50 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X286 GND word49 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X287 Y3 word34 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X288 GND word21 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X289 Y4 word110 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X290 GND word101 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X291 Y0 word94 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X292 GND word119 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X293 Y6 word16 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X294 Y7 word44 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X295 GND word121 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X296 Y2 word114 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X297 GND word103 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X298 GND word87 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X299 Y0 word56 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X300 GND word43 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X301 GND word45 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X302 GND word23 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X303 GND word25 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X304 Y3 word28 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X305 GND word27 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X306 Y3 word112 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X307 Y6 word94 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X308 GND word101 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X309 GND word55 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X310 Y3 word92 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X311 Y1 word116 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X312 Y7 word110 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X313 Y1 word98 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X314 GND word69 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X315 Y3 word54 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X316 Y4 word52 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X317 GND word65 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X318 GND word87 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X319 Y5 word20 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X320 Y1 word36 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X321 Y1 word18 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X322 Y4 word112 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X323 Y0 word114 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X324 Y7 word46 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X325 Y4 word92 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X326 GND word107 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X327 Y2 word60 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X328 GND word45 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X329 Y2 word42 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X330 GND word47 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X331 GND word27 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X332 GND word29 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X333 Y6 word114 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X334 GND word87 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X335 Y6 word24 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X336 Y7 word112 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X337 GND word21 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X338 GND word107 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X339 GND word111 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X340 Y5 word40 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X341 Y7 word92 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X342 GND word67 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X343 GND word51 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X344 Y3 word36 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X345 Y1 word38 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X346 Y3 word74 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X347 Y3 word18 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X348 Y7 word48 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X349 Y2 word16 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X350 Y2 word62 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X351 Y4 word60 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X352 Y4 word42 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X353 GND word47 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X354 GND word31 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X355 Y0 word58 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X356 Y6 word116 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X357 Y1 word44 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X358 GND word111 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X359 Y6 word26 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X360 GND word85 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X361 Y2 word124 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X362 GND word115 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X363 Y0 word20 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X364 Y3 word76 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X365 GND word55 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X366 GND word53 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X367 Y3 word38 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X368 Y5 word22 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X369 GND word107 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X370 GND word19 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X371 GND word111 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X372 Y1 word126 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X373 Y4 word16 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X374 GND word17 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X375 Y4 word62 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X376 GND word29 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X377 Y3 word44 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X378 Y1 word46 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X379 Y0 word124 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X380 Y4 word76 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X381 GND word71 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X382 Y0 word40 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X383 GND word117 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X384 Y2 word24 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X385 GND word111 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X386 Y2 word70 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X387 GND word113 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X388 GND word55 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X389 GND word39 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X390 GND word37 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X391 Y3 word122 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X392 Y5 word78 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X393 GND word31 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X394 Y7 word120 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X395 GND word71 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X396 Y1 word108 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X397 GND word117 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X398 Y1 word66 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X399 Y3 word84 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X400 GND word61 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X401 Y3 word46 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X402 Y1 word48 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X403 Y5 word30 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X404 GND word115 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X405 GND word113 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X406 GND word85 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X407 Y4 word24 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X408 GND word25 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X409 Y6 word28 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X410 Y2 word26 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X411 Y0 word22 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X412 Y0 word68 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X413 GND word57 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X414 GND word37 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X415 Y4 word84 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X416 Y3 word78 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X417 GND word71 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X418 GND word21 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X419 GND word113 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X420 GND word95 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X421 GND word79 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X422 GND word77 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X423 GND word33 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X424 GND word35 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X425 GND word17 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X426 GND word19 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X427 Y3 word66 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X428 GND word63 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X429 Y3 word48 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X430 GND word117 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X431 GND word75 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X432 Y1 word90 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X433 GND word45 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X434 Y7 word84 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X435 Y4 word26 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X436 GND word27 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X437 Y5 word86 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X438 GND word39 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X439 GND word79 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X440 GND word113 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X441 GND word125 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X442 GND word57 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X443 Y1 word56 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X444 GND word23 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X445 Y6 word108 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X446 Y7 word20 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X447 Y2 word90 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X448 GND word81 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X449 GND word17 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X450 Y6 word18 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X451 GND word19 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X452 Y2 word34 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X453 Y0 word30 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X454 GND word123 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X455 Y5 word52 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X456 GND word49 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X457 GND word95 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X458 GND word65 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X459 Y3 word86 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X460 GND word79 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X461 GND word125 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X462 Y7 word104 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X463 GND word29 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X464 GND word47 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X465 Y5 word88 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X466 GND word59 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X467 GND word81 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X468 Y1 word72 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X469 GND word41 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X470 GND word25 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X471 Y2 word28 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X472 Y0 word90 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X473 Y3 word56 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X474 GND word43 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X475 GND word79 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X476 GND word123 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X477 GND word95 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X478 GND word83 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X479 Y6 word38 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X480 Y2 word54 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X481 Y4 word34 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X482 Y5 word94 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X483 GND word127 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X484 Y0 word50 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X485 Y2 word72 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X486 GND word69 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X487 GND word21 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X488 Y6 word90 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X489 Y3 word88 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X490 GND word67 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X491 GND word81 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X492 GND word31 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X493 GND word123 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X494 GND word89 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X495 Y7 word86 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X496 GND word45 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X497 GND word83 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X498 Y4 word28 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X499 GND word25 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X500 GND word27 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X501 Y5 word60 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X502 GND word23 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X503 VDD GND Y6 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X504 Y3 word94 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X505 Y1 word58 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X506 Y4 word88 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X507 Y0 word72 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X508 Y7 word22 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X509 Y5 word114 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X510 Y4 word54 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X511 GND word89 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X512 Y1 word80 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X513 Y0 word52 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X514 GND word49 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X515 Y2 word36 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X516 Y1 word20 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X517 GND word21 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X518 Y2 word18 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X519 GND word105 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X520 GND word83 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X521 GND word109 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X522 GND word91 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X523 Y6 word46 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X524 Y7 word88 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X525 GND word47 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X526 GND word27 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X527 GND word87 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X528 Y5 word16 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X529 GND word43 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X530 Y2 word80 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X531 GND word29 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X532 GND word105 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X533 Y3 word58 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X534 GND word89 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X535 Y7 word94 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X536 GND word69 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X537 GND word91 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X538 Y1 word82 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X539 Y4 word36 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X540 GND word37 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X541 Y2 word38 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X542 Y1 word40 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X543 Y4 word18 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X544 Y3 word20 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X545 Y4 word114 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X546 GND word89 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X547 GND word53 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X548 Y0 word80 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X549 GND word105 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X550 Y7 word30 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X551 Y6 word48 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X552 Y2 word100 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X553 Y0 word60 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X554 Y2 word82 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X555 Y0 word42 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X556 Y2 word44 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X557 GND word73 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X558 GND word29 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X559 GND word31 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X560 Y3 word116 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X561 Y3 word98 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X562 GND word91 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X563 Y6 word80 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X564 GND word41 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X565 GND word87 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X566 Y7 word114 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X567 Y1 word102 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X568 GND word57 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X569 GND word55 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X570 Y4 word38 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X571 Y3 word40 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X572 Y5 word24 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X573 GND word51 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X574 GND word109 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X575 GND word73 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X576 Y5 word70 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X577 Y1 word22 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X578 Y4 word116 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X579 GND word91 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X580 Y0 word100 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X581 Y1 word68 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X582 Y0 word82 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X583 GND word19 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X584 Y7 word50 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X585 Y5 word124 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X586 Y0 word16 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X587 Y2 word102 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X588 GND word93 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X589 Y0 word62 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X590 Y4 word44 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X591 Y2 word46 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X592 GND word87 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X593 GND word31 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X594 GND word33 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X595 GND word61 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X596 VDD GND Y4 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X597 Y7 word116 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X598 GND word73 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X599 GND word115 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X600 Y6 word56 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X601 GND word23 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X602 GND word93 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X603 Y5 word26 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X604 GND word53 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X605 GND word37 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X606 GND word39 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X607 Y3 word22 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X608 Y0 word102 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X609 Y3 word68 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
*.ends

