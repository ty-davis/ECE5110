magic
tech sky130A
magscale 1 2
timestamp 1744838505
<< nwell >>
rect -54 -17586 1946 -17176
<< nmos >>
rect 978 -17986 1080 -17952
rect 1476 -17986 1578 -17952
rect 1476 -18128 1578 -18094
<< pmos >>
rect -18 -17450 84 -17416
rect 314 -17450 416 -17416
rect 480 -17450 582 -17416
rect 812 -17450 914 -17416
rect 978 -17450 1080 -17416
rect 1310 -17450 1412 -17416
rect 1476 -17450 1578 -17416
rect 1808 -17450 1910 -17416
<< ndiff >>
rect 978 -17880 1080 -17864
rect 978 -17914 1012 -17880
rect 1046 -17914 1080 -17880
rect 978 -17952 1080 -17914
rect 1476 -17880 1578 -17864
rect 1476 -17914 1510 -17880
rect 1544 -17914 1578 -17880
rect 1476 -17952 1578 -17914
rect 978 -18006 1080 -17986
rect 1476 -18006 1578 -17986
rect 978 -18022 1228 -18006
rect 978 -18056 1178 -18022
rect 1212 -18056 1228 -18022
rect 978 -18072 1228 -18056
rect 1476 -18022 1726 -18006
rect 1476 -18056 1676 -18022
rect 1710 -18056 1726 -18022
rect 1476 -18072 1726 -18056
rect 1476 -18094 1578 -18072
rect 1476 -18164 1578 -18128
rect 1476 -18198 1510 -18164
rect 1544 -18198 1578 -18164
rect 1476 -18214 1578 -18198
<< pdiff >>
rect -18 -17340 84 -17322
rect -18 -17394 -2 -17340
rect 66 -17394 84 -17340
rect -18 -17416 84 -17394
rect 314 -17340 416 -17322
rect 314 -17394 330 -17340
rect 398 -17394 416 -17340
rect 314 -17416 416 -17394
rect 480 -17340 582 -17322
rect 480 -17394 496 -17340
rect 564 -17394 582 -17340
rect 480 -17416 582 -17394
rect 812 -17340 914 -17322
rect 812 -17394 828 -17340
rect 896 -17394 914 -17340
rect 812 -17416 914 -17394
rect 978 -17340 1080 -17322
rect 978 -17394 994 -17340
rect 1062 -17394 1080 -17340
rect 978 -17416 1080 -17394
rect 1310 -17340 1412 -17322
rect 1310 -17394 1326 -17340
rect 1394 -17394 1412 -17340
rect 1310 -17416 1412 -17394
rect 1476 -17340 1578 -17322
rect 1476 -17394 1492 -17340
rect 1560 -17394 1578 -17340
rect 1476 -17416 1578 -17394
rect 1808 -17340 1910 -17322
rect 1808 -17394 1824 -17340
rect 1892 -17394 1910 -17340
rect 1808 -17416 1910 -17394
rect -18 -17472 84 -17450
rect -18 -17506 16 -17472
rect 50 -17506 84 -17472
rect -18 -17522 84 -17506
rect 314 -17472 416 -17450
rect 314 -17506 348 -17472
rect 382 -17506 416 -17472
rect 314 -17522 416 -17506
rect 480 -17472 582 -17450
rect 480 -17506 514 -17472
rect 548 -17506 582 -17472
rect 480 -17522 582 -17506
rect 812 -17472 914 -17450
rect 812 -17506 846 -17472
rect 880 -17506 914 -17472
rect 812 -17522 914 -17506
rect 978 -17472 1080 -17450
rect 978 -17506 1012 -17472
rect 1046 -17506 1080 -17472
rect 978 -17522 1080 -17506
rect 1310 -17472 1412 -17450
rect 1310 -17506 1344 -17472
rect 1378 -17506 1412 -17472
rect 1310 -17522 1412 -17506
rect 1476 -17472 1578 -17450
rect 1476 -17506 1510 -17472
rect 1544 -17506 1578 -17472
rect 1476 -17522 1578 -17506
rect 1808 -17472 1910 -17450
rect 1808 -17506 1842 -17472
rect 1876 -17506 1910 -17472
rect 1808 -17522 1910 -17506
<< ndiffc >>
rect 1012 -17914 1046 -17880
rect 1510 -17914 1544 -17880
rect 1178 -18056 1212 -18022
rect 1676 -18056 1710 -18022
rect 1510 -18198 1544 -18164
<< pdiffc >>
rect -2 -17394 66 -17340
rect 330 -17394 398 -17340
rect 496 -17394 564 -17340
rect 828 -17394 896 -17340
rect 994 -17394 1062 -17340
rect 1326 -17394 1394 -17340
rect 1492 -17394 1560 -17340
rect 1824 -17394 1892 -17340
rect 16 -17506 50 -17472
rect 348 -17506 382 -17472
rect 514 -17506 548 -17472
rect 846 -17506 880 -17472
rect 1012 -17506 1046 -17472
rect 1344 -17506 1378 -17472
rect 1510 -17506 1544 -17472
rect 1842 -17506 1876 -17472
<< psubdiff >>
rect -54 -17792 -30 -17736
rect 1702 -17792 1726 -17736
<< nsubdiff >>
rect -18 -17268 6 -17212
rect 1886 -17268 1910 -17212
<< psubdiffcont >>
rect -30 -17792 1702 -17736
<< nsubdiffcont >>
rect 6 -17268 1886 -17212
<< poly >>
rect -120 -17416 -54 -17400
rect -120 -17450 -104 -17416
rect -70 -17450 -18 -17416
rect 84 -17450 314 -17416
rect 416 -17450 480 -17416
rect 582 -17450 812 -17416
rect 914 -17450 978 -17416
rect 1080 -17450 1310 -17416
rect 1412 -17450 1476 -17416
rect 1578 -17450 1808 -17416
rect 1910 -17450 1936 -17416
rect -120 -17466 -54 -17450
rect -118 -17952 -52 -17936
rect -118 -17986 -102 -17952
rect -68 -17986 978 -17952
rect 1080 -17986 1476 -17952
rect 1578 -17986 1992 -17952
rect -118 -18002 -52 -17986
rect -118 -18094 -52 -18078
rect -118 -18128 -102 -18094
rect -68 -18128 1476 -18094
rect 1578 -18128 1992 -18094
rect -118 -18144 -52 -18128
<< polycont >>
rect -104 -17450 -70 -17416
rect -102 -17986 -68 -17952
rect -102 -18128 -68 -18094
<< locali >>
rect -50 -17212 1942 -17192
rect -50 -17268 6 -17212
rect 1886 -17268 1942 -17212
rect -50 -17288 1942 -17268
rect -18 -17340 84 -17288
rect -18 -17394 -2 -17340
rect 66 -17394 84 -17340
rect -120 -17416 -54 -17400
rect -18 -17410 84 -17394
rect 314 -17340 416 -17288
rect 314 -17394 330 -17340
rect 398 -17394 416 -17340
rect 314 -17410 416 -17394
rect 480 -17340 582 -17288
rect 480 -17394 496 -17340
rect 564 -17394 582 -17340
rect 480 -17410 582 -17394
rect 812 -17340 914 -17288
rect 812 -17394 828 -17340
rect 896 -17394 914 -17340
rect 812 -17410 914 -17394
rect 978 -17340 1080 -17288
rect 978 -17394 994 -17340
rect 1062 -17394 1080 -17340
rect 978 -17410 1080 -17394
rect 1310 -17340 1412 -17288
rect 1310 -17394 1326 -17340
rect 1394 -17394 1412 -17340
rect 1310 -17410 1412 -17394
rect 1476 -17340 1578 -17288
rect 1476 -17394 1492 -17340
rect 1560 -17394 1578 -17340
rect 1476 -17410 1578 -17394
rect 1808 -17340 1910 -17288
rect 1808 -17394 1824 -17340
rect 1892 -17394 1910 -17340
rect 1808 -17410 1910 -17394
rect -120 -17450 -104 -17416
rect -70 -17450 -54 -17416
rect -120 -17716 -54 -17450
rect 0 -17472 66 -17456
rect 0 -17506 16 -17472
rect 50 -17506 66 -17472
rect 0 -17522 66 -17506
rect 332 -17472 398 -17456
rect 332 -17506 348 -17472
rect 382 -17506 398 -17472
rect 332 -17522 398 -17506
rect 498 -17472 564 -17456
rect 498 -17506 514 -17472
rect 548 -17506 564 -17472
rect 498 -17522 564 -17506
rect 830 -17472 896 -17456
rect 830 -17506 846 -17472
rect 880 -17506 896 -17472
rect 830 -17522 896 -17506
rect 996 -17472 1062 -17456
rect 996 -17506 1012 -17472
rect 1046 -17506 1062 -17472
rect 996 -17522 1062 -17506
rect 1328 -17472 1394 -17456
rect 1328 -17506 1344 -17472
rect 1378 -17506 1394 -17472
rect 1328 -17522 1394 -17506
rect 1494 -17472 1560 -17456
rect 1494 -17506 1510 -17472
rect 1544 -17506 1560 -17472
rect 1494 -17522 1560 -17506
rect 1826 -17472 1892 -17456
rect 1826 -17506 1842 -17472
rect 1876 -17506 1892 -17472
rect 1826 -17522 1892 -17506
rect -120 -17736 1726 -17716
rect -120 -17792 -30 -17736
rect 1702 -17792 1726 -17736
rect -120 -17812 1726 -17792
rect 166 -17834 234 -17812
rect 662 -17834 732 -17812
rect 1162 -17834 1230 -17812
rect 0 -17862 66 -17846
rect 0 -17896 16 -17862
rect 50 -17896 66 -17862
rect -118 -17952 -52 -17936
rect -118 -17986 -102 -17952
rect -68 -17986 -52 -17952
rect -118 -18002 -52 -17986
rect -118 -18094 -52 -18078
rect -118 -18128 -102 -18094
rect -68 -18128 -52 -18094
rect -118 -18144 -52 -18128
rect 0 -18236 66 -17896
rect 166 -17883 233 -17834
rect 332 -17862 398 -17846
rect 166 -18236 232 -17883
rect 332 -17896 348 -17862
rect 382 -17896 398 -17862
rect 332 -18236 398 -17896
rect 498 -17862 564 -17846
rect 498 -17896 514 -17862
rect 548 -17896 564 -17862
rect 498 -18236 564 -17896
rect 663 -17909 730 -17834
rect 664 -18236 730 -17909
rect 830 -17862 896 -17846
rect 830 -17896 846 -17862
rect 880 -17896 896 -17862
rect 830 -18236 896 -17896
rect 996 -17862 1062 -17846
rect 996 -17914 1012 -17862
rect 1046 -17914 1062 -17862
rect 996 -18236 1062 -17914
rect 1162 -17885 1229 -17834
rect 1328 -17862 1394 -17846
rect 1162 -18022 1228 -17885
rect 1162 -18056 1178 -18022
rect 1212 -18056 1228 -18022
rect 1162 -18236 1228 -18056
rect 1328 -17896 1344 -17862
rect 1378 -17896 1394 -17862
rect 1328 -18236 1394 -17896
rect 1494 -17862 1560 -17846
rect 1494 -17914 1510 -17862
rect 1544 -17914 1560 -17862
rect 1494 -18164 1560 -17914
rect 1494 -18198 1510 -18164
rect 1544 -18198 1560 -18164
rect 1494 -18236 1560 -18198
rect 1660 -18022 1726 -17812
rect 1660 -18056 1676 -18022
rect 1710 -18056 1726 -18022
rect 1660 -18236 1726 -18056
rect 1826 -17862 1892 -17846
rect 1826 -17896 1842 -17862
rect 1876 -17896 1892 -17862
rect 1826 -18236 1892 -17896
<< viali >>
rect 16 -17506 50 -17472
rect 348 -17506 382 -17472
rect 514 -17506 548 -17472
rect 846 -17506 880 -17472
rect 1012 -17506 1046 -17472
rect 1344 -17506 1378 -17472
rect 1510 -17506 1544 -17472
rect 1842 -17506 1876 -17472
rect 16 -17896 50 -17862
rect 348 -17896 382 -17862
rect 514 -17896 548 -17862
rect 846 -17896 880 -17862
rect 1012 -17880 1046 -17862
rect 1012 -17896 1046 -17880
rect 1344 -17896 1378 -17862
rect 1510 -17880 1544 -17862
rect 1510 -17896 1544 -17880
rect 1842 -17896 1876 -17862
<< metal1 >>
rect 0 -17472 66 -17456
rect 0 -17506 16 -17472
rect 50 -17506 66 -17472
rect 0 -17862 66 -17506
rect 0 -17896 16 -17862
rect 50 -17896 66 -17862
rect 0 -17912 66 -17896
rect 332 -17472 398 -17456
rect 332 -17506 348 -17472
rect 382 -17506 398 -17472
rect 332 -17862 398 -17506
rect 332 -17896 348 -17862
rect 382 -17896 398 -17862
rect 332 -17912 398 -17896
rect 498 -17472 564 -17456
rect 498 -17506 514 -17472
rect 548 -17506 564 -17472
rect 498 -17862 564 -17506
rect 498 -17896 514 -17862
rect 548 -17896 564 -17862
rect 498 -17912 564 -17896
rect 830 -17472 896 -17456
rect 830 -17506 846 -17472
rect 880 -17506 896 -17472
rect 830 -17862 896 -17506
rect 830 -17896 846 -17862
rect 880 -17896 896 -17862
rect 830 -17912 896 -17896
rect 996 -17472 1062 -17456
rect 996 -17506 1012 -17472
rect 1046 -17506 1062 -17472
rect 996 -17862 1062 -17506
rect 996 -17896 1012 -17862
rect 1046 -17896 1062 -17862
rect 996 -17912 1062 -17896
rect 1328 -17472 1394 -17456
rect 1328 -17506 1344 -17472
rect 1378 -17506 1394 -17472
rect 1328 -17862 1394 -17506
rect 1328 -17896 1344 -17862
rect 1378 -17896 1394 -17862
rect 1328 -17912 1394 -17896
rect 1494 -17472 1560 -17456
rect 1494 -17506 1510 -17472
rect 1544 -17506 1560 -17472
rect 1494 -17862 1560 -17506
rect 1494 -17896 1510 -17862
rect 1544 -17896 1560 -17862
rect 1494 -17912 1560 -17896
rect 1826 -17472 1892 -17456
rect 1826 -17506 1842 -17472
rect 1876 -17506 1892 -17472
rect 1826 -17862 1892 -17506
rect 1826 -17896 1842 -17862
rect 1876 -17896 1892 -17862
rect 1826 -17912 1892 -17896
<< labels >>
flabel locali -118 -18002 -52 -17936 0 FreeSerif 160 0 0 0 word126
port 32 nsew
flabel locali -118 -18144 -52 -18078 0 FreeSerif 160 0 0 0 word127
port 35 nsew
flabel locali 332 -18236 398 -18170 0 FreeSerif 160 0 0 0 Y6
port 38 nsew
flabel locali 0 -18236 66 -18170 0 FreeSerif 160 0 0 0 Y7
port 37 nsew
flabel locali 498 -18236 564 -18170 0 FreeSerif 160 0 0 0 Y5
port 39 nsew
flabel locali 830 -18236 896 -18170 0 FreeSerif 160 0 0 0 Y4
port 40 nsew
flabel locali 996 -18236 1062 -18170 0 FreeSerif 160 0 0 0 Y3
port 41 nsew
flabel locali 1328 -18236 1394 -18170 0 FreeSerif 160 0 0 0 Y2
port 42 nsew
flabel locali 1494 -18236 1560 -18170 0 FreeSerif 160 0 0 0 Y1
port 43 nsew
flabel locali 1826 -18236 1892 -18170 0 FreeSerif 160 0 0 0 Y0
port 44 nsew
flabel locali 132 -17812 278 -17716 0 FreeSerif 160 0 0 0 GND!
port 0 nsew
flabel locali -50 -17288 1942 -17192 0 FreeSerif 160 0 0 0 VDD!
port 10 nsew
<< end >>
