magic
tech sky130A
timestamp 1741888123
<< error_p >>
rect 185 315 208 415
rect 185 65 208 115
rect 313 -130 325 -118
rect 326 -130 343 -112
rect 308 -142 343 -130
rect 308 -146 325 -142
rect 326 -146 343 -142
rect 308 -158 343 -146
rect 313 -170 325 -158
rect 326 -176 343 -158
rect 315 -562 327 -550
rect 327 -574 339 -562
rect 327 -590 339 -578
rect 315 -602 327 -590
<< nwell >>
rect -2 197 796 488
rect -2 -403 326 -112
<< nmos >>
rect 72 65 87 115
rect 126 65 141 115
rect 210 65 225 115
rect 264 65 279 115
rect 438 65 453 115
rect 492 65 507 115
rect 613 65 628 115
rect 667 65 682 115
rect 72 -535 87 -485
rect 126 -535 141 -485
rect 179 -535 194 -485
rect 233 -535 248 -485
<< pmos >>
rect 72 315 87 415
rect 126 315 141 415
rect 210 315 225 415
rect 264 315 279 415
rect 438 315 453 415
rect 492 315 507 415
rect 613 315 628 415
rect 667 315 682 415
rect 72 -285 87 -185
rect 126 -285 141 -185
rect 179 -285 194 -185
rect 233 -285 248 -185
<< ndiff >>
rect 36 107 72 115
rect 36 73 44 107
rect 61 73 72 107
rect 36 65 72 73
rect 87 107 126 115
rect 87 73 98 107
rect 115 73 126 107
rect 87 65 126 73
rect 141 107 177 115
rect 141 73 152 107
rect 169 73 177 107
rect 141 65 177 73
rect 208 65 210 115
rect 225 107 264 115
rect 225 73 236 107
rect 253 73 264 107
rect 225 65 264 73
rect 279 107 315 115
rect 279 73 290 107
rect 307 73 315 107
rect 279 65 315 73
rect 402 107 438 115
rect 402 73 410 107
rect 427 73 438 107
rect 402 65 438 73
rect 453 107 492 115
rect 453 73 464 107
rect 481 73 492 107
rect 453 65 492 73
rect 507 107 543 115
rect 507 73 518 107
rect 535 73 543 107
rect 507 65 543 73
rect 577 107 613 115
rect 577 73 585 107
rect 602 73 613 107
rect 577 65 613 73
rect 628 107 667 115
rect 628 73 639 107
rect 656 73 667 107
rect 628 65 667 73
rect 682 107 718 115
rect 682 73 693 107
rect 710 73 718 107
rect 682 65 718 73
rect 36 -493 72 -485
rect 36 -527 44 -493
rect 61 -527 72 -493
rect 36 -535 72 -527
rect 87 -493 126 -485
rect 87 -527 98 -493
rect 115 -527 126 -493
rect 87 -535 126 -527
rect 141 -493 179 -485
rect 141 -527 152 -493
rect 169 -527 179 -493
rect 141 -535 179 -527
rect 194 -493 233 -485
rect 194 -527 205 -493
rect 222 -527 233 -493
rect 194 -535 233 -527
rect 248 -493 284 -485
rect 248 -527 259 -493
rect 276 -527 284 -493
rect 248 -535 284 -527
<< pdiff >>
rect 36 407 72 415
rect 36 323 44 407
rect 61 323 72 407
rect 36 315 72 323
rect 87 407 126 415
rect 87 323 98 407
rect 115 323 126 407
rect 87 315 126 323
rect 141 407 177 415
rect 141 323 152 407
rect 169 323 177 407
rect 141 315 177 323
rect 208 315 210 415
rect 225 407 264 415
rect 225 323 236 407
rect 253 323 264 407
rect 225 315 264 323
rect 279 407 315 415
rect 279 323 290 407
rect 307 323 315 407
rect 279 315 315 323
rect 402 407 438 415
rect 402 323 410 407
rect 427 323 438 407
rect 402 315 438 323
rect 453 407 492 415
rect 453 323 464 407
rect 481 323 492 407
rect 453 315 492 323
rect 507 407 543 415
rect 507 323 518 407
rect 535 323 543 407
rect 507 315 543 323
rect 577 407 613 415
rect 577 323 585 407
rect 602 323 613 407
rect 577 315 613 323
rect 628 407 667 415
rect 628 323 639 407
rect 656 323 667 407
rect 628 315 667 323
rect 682 407 718 415
rect 682 323 693 407
rect 710 323 718 407
rect 682 315 718 323
rect 36 -193 72 -185
rect 36 -277 44 -193
rect 61 -277 72 -193
rect 36 -285 72 -277
rect 87 -193 126 -185
rect 87 -277 98 -193
rect 115 -277 126 -193
rect 87 -285 126 -277
rect 141 -193 179 -185
rect 141 -277 152 -193
rect 169 -277 179 -193
rect 141 -285 179 -277
rect 194 -193 233 -185
rect 194 -277 205 -193
rect 222 -277 233 -193
rect 194 -285 233 -277
rect 248 -193 284 -185
rect 248 -277 259 -193
rect 276 -277 284 -193
rect 248 -285 284 -277
<< ndiffc >>
rect 44 73 61 107
rect 98 73 115 107
rect 152 73 169 107
rect 236 73 253 107
rect 290 73 307 107
rect 410 73 427 107
rect 464 73 481 107
rect 518 73 535 107
rect 585 73 602 107
rect 639 73 656 107
rect 693 73 710 107
rect 44 -527 61 -493
rect 98 -527 115 -493
rect 152 -527 169 -493
rect 205 -527 222 -493
rect 259 -527 276 -493
<< pdiffc >>
rect 44 323 61 407
rect 98 323 115 407
rect 152 323 169 407
rect 236 323 253 407
rect 290 323 307 407
rect 410 323 427 407
rect 464 323 481 407
rect 518 323 535 407
rect 585 323 602 407
rect 639 323 656 407
rect 693 323 710 407
rect 44 -277 61 -193
rect 98 -277 115 -193
rect 152 -277 169 -193
rect 205 -277 222 -193
rect 259 -277 276 -193
<< psubdiff >>
rect 0 10 12 38
rect 782 10 794 38
rect 0 -590 12 -562
<< nsubdiff >>
rect 16 442 28 470
rect 766 442 778 470
rect 16 -158 28 -130
<< psubdiffcont >>
rect 12 10 782 38
rect 12 -590 327 -562
<< nsubdiffcont >>
rect 28 442 766 470
rect 28 -158 325 -130
<< poly >>
rect 72 415 87 428
rect 126 415 141 428
rect 210 415 225 428
rect 264 415 279 428
rect 438 415 453 428
rect 492 415 507 428
rect 613 415 628 428
rect 667 415 682 428
rect 72 224 87 315
rect 126 282 141 315
rect 126 274 159 282
rect 126 257 134 274
rect 151 257 159 274
rect 126 249 159 257
rect 72 207 141 224
rect 115 199 141 207
rect 42 175 75 183
rect 42 158 50 175
rect 67 158 75 175
rect 126 182 141 199
rect 210 223 225 315
rect 264 278 279 315
rect 438 295 453 315
rect 420 287 453 295
rect 247 270 280 278
rect 247 253 255 270
rect 272 263 280 270
rect 420 270 428 287
rect 445 270 453 287
rect 272 253 316 263
rect 420 262 453 270
rect 247 245 316 253
rect 210 215 243 223
rect 210 198 218 215
rect 235 198 243 215
rect 210 190 243 198
rect 126 174 159 182
rect 42 150 87 158
rect 57 139 87 150
rect 72 115 87 139
rect 126 157 134 174
rect 151 157 159 174
rect 126 149 159 157
rect 126 115 141 149
rect 210 115 225 190
rect 297 151 316 245
rect 492 228 507 315
rect 613 276 628 315
rect 613 268 646 276
rect 613 259 621 268
rect 418 216 507 228
rect 405 213 507 216
rect 578 251 621 259
rect 638 251 646 268
rect 578 243 646 251
rect 405 208 438 213
rect 405 191 413 208
rect 430 191 438 208
rect 405 183 438 191
rect 264 132 316 151
rect 418 150 438 183
rect 492 184 525 192
rect 492 167 500 184
rect 517 167 525 184
rect 492 159 525 167
rect 418 135 453 150
rect 264 115 279 132
rect 438 115 453 135
rect 492 115 507 159
rect 578 144 596 243
rect 667 218 682 315
rect 634 210 682 218
rect 634 193 642 210
rect 659 193 682 210
rect 634 185 682 193
rect 578 129 628 144
rect 613 115 628 129
rect 667 115 682 185
rect 72 52 87 65
rect 126 52 141 65
rect 210 52 225 65
rect 264 52 279 65
rect 438 52 453 65
rect 492 52 507 65
rect 613 52 628 65
rect 667 52 682 65
rect 72 -185 87 -172
rect 126 -185 141 -172
rect 179 -185 194 -172
rect 233 -185 248 -172
rect 72 -305 87 -285
rect 72 -313 105 -305
rect 72 -330 80 -313
rect 97 -330 105 -313
rect 72 -338 105 -330
rect 72 -399 87 -338
rect 126 -345 141 -285
rect 125 -353 158 -345
rect 125 -370 133 -353
rect 150 -370 158 -353
rect 125 -378 158 -370
rect 72 -414 141 -399
rect 72 -443 105 -435
rect 72 -460 80 -443
rect 97 -460 105 -443
rect 72 -468 105 -460
rect 72 -485 87 -468
rect 126 -485 141 -414
rect 179 -435 194 -285
rect 233 -381 248 -285
rect 215 -389 248 -381
rect 215 -406 223 -389
rect 240 -406 248 -389
rect 215 -414 248 -406
rect 179 -443 212 -435
rect 179 -460 187 -443
rect 204 -460 212 -443
rect 179 -468 212 -460
rect 179 -485 194 -468
rect 233 -485 248 -414
rect 72 -548 87 -535
rect 126 -548 141 -535
rect 179 -548 194 -535
rect 233 -548 248 -535
<< polycont >>
rect 134 257 151 274
rect 50 158 67 175
rect 255 253 272 270
rect 428 270 445 287
rect 218 198 235 215
rect 134 157 151 174
rect 621 251 638 268
rect 413 191 430 208
rect 500 167 517 184
rect 642 193 659 210
rect 80 -330 97 -313
rect 133 -370 150 -353
rect 80 -460 97 -443
rect 223 -406 240 -389
rect 187 -460 204 -443
<< locali >>
rect 0 470 794 480
rect 0 442 28 470
rect 766 442 794 470
rect 0 432 794 442
rect 36 407 69 415
rect 36 323 44 407
rect 61 323 69 407
rect 36 315 69 323
rect 90 407 123 415
rect 90 323 98 407
rect 115 323 123 407
rect 90 315 123 323
rect 144 407 177 415
rect 144 323 152 407
rect 169 323 177 407
rect 144 316 177 323
rect 228 407 261 432
rect 228 323 236 407
rect 253 323 261 407
rect 36 272 58 315
rect 7 264 58 272
rect 7 247 15 264
rect 32 256 58 264
rect 32 255 54 256
rect 32 247 40 255
rect 7 239 40 247
rect 8 133 25 239
rect 92 232 109 315
rect 144 299 193 316
rect 228 315 261 323
rect 282 407 315 415
rect 282 323 290 407
rect 307 323 315 407
rect 402 407 435 415
rect 402 332 410 407
rect 282 315 315 323
rect 126 274 159 282
rect 126 257 134 274
rect 151 257 159 274
rect 126 249 159 257
rect 92 224 128 232
rect 42 209 75 216
rect 42 192 50 209
rect 67 192 75 209
rect 42 175 75 192
rect 42 158 50 175
rect 67 158 75 175
rect 42 150 75 158
rect 92 207 103 224
rect 120 207 128 224
rect 92 199 128 207
rect 8 115 69 133
rect 92 119 109 199
rect 126 174 159 182
rect 126 157 134 174
rect 151 157 159 174
rect 126 149 159 157
rect 176 132 193 299
rect 247 270 280 278
rect 247 253 255 270
rect 272 253 280 270
rect 247 245 280 253
rect 210 215 243 223
rect 210 198 218 215
rect 235 207 243 215
rect 297 207 315 315
rect 385 323 410 332
rect 427 323 435 407
rect 385 315 435 323
rect 456 407 489 415
rect 456 323 464 407
rect 481 323 489 407
rect 456 315 489 323
rect 385 267 402 315
rect 235 198 315 207
rect 210 190 315 198
rect 36 107 69 115
rect 36 73 44 107
rect 61 73 69 107
rect 36 65 69 73
rect 90 107 123 119
rect 90 73 98 107
rect 115 73 123 107
rect 90 65 123 73
rect 144 115 193 132
rect 282 182 315 190
rect 369 259 402 267
rect 420 287 453 295
rect 420 270 428 287
rect 445 270 453 287
rect 420 262 453 270
rect 369 242 377 259
rect 394 242 402 259
rect 472 261 489 315
rect 510 407 543 415
rect 510 323 518 407
rect 535 323 543 407
rect 510 316 543 323
rect 577 407 610 415
rect 577 323 585 407
rect 602 323 610 407
rect 510 299 560 316
rect 472 253 505 261
rect 472 245 480 253
rect 369 234 402 242
rect 456 236 480 245
rect 497 236 505 253
rect 282 115 300 182
rect 369 133 386 234
rect 456 228 505 236
rect 405 208 438 216
rect 405 191 413 208
rect 430 191 438 208
rect 405 175 438 191
rect 405 158 413 175
rect 430 158 438 175
rect 405 150 438 158
rect 369 115 435 133
rect 144 107 177 115
rect 144 73 152 107
rect 169 73 177 107
rect 144 65 177 73
rect 228 107 261 115
rect 228 73 236 107
rect 253 73 261 107
rect 228 48 261 73
rect 282 107 315 115
rect 282 73 290 107
rect 307 73 315 107
rect 282 65 315 73
rect 402 107 435 115
rect 402 73 410 107
rect 427 73 435 107
rect 402 65 435 73
rect 456 115 473 228
rect 492 184 525 192
rect 492 167 500 184
rect 517 167 525 184
rect 492 159 525 167
rect 542 165 560 299
rect 577 315 610 323
rect 631 407 664 432
rect 631 323 639 407
rect 656 323 664 407
rect 631 315 664 323
rect 685 407 718 415
rect 685 323 693 407
rect 710 323 718 407
rect 577 209 594 315
rect 613 268 646 276
rect 613 251 621 268
rect 638 251 646 268
rect 613 243 646 251
rect 634 210 667 218
rect 577 203 610 209
rect 634 203 642 210
rect 577 193 642 203
rect 659 193 667 210
rect 577 192 667 193
rect 593 185 667 192
rect 542 157 575 165
rect 542 140 550 157
rect 567 140 575 157
rect 542 132 575 140
rect 510 115 560 132
rect 593 115 610 185
rect 685 157 718 323
rect 685 140 693 157
rect 710 140 718 157
rect 456 107 489 115
rect 456 73 464 107
rect 481 73 489 107
rect 456 65 489 73
rect 510 107 543 115
rect 510 73 518 107
rect 535 73 543 107
rect 510 65 543 73
rect 577 107 610 115
rect 577 73 585 107
rect 602 73 610 107
rect 577 65 610 73
rect 631 107 664 115
rect 631 73 639 107
rect 656 73 664 107
rect 631 48 664 73
rect 685 107 718 140
rect 685 73 693 107
rect 710 73 718 107
rect 685 65 718 73
rect 0 38 794 48
rect 0 10 12 38
rect 782 10 794 38
rect 0 0 794 10
rect 0 -130 325 -120
rect 0 -158 28 -130
rect 0 -168 325 -158
rect 36 -193 69 -185
rect 36 -277 44 -193
rect 61 -277 69 -193
rect 36 -285 69 -277
rect 90 -193 123 -185
rect 90 -277 98 -193
rect 115 -277 123 -193
rect 90 -285 123 -277
rect 144 -193 177 -185
rect 144 -277 152 -193
rect 169 -277 177 -193
rect 144 -285 177 -277
rect 197 -193 230 -168
rect 197 -277 205 -193
rect 222 -277 230 -193
rect 197 -285 230 -277
rect 251 -193 284 -185
rect 251 -277 259 -193
rect 276 -277 284 -193
rect 251 -285 284 -277
rect 36 -485 53 -285
rect 160 -302 177 -285
rect 72 -313 105 -305
rect 72 -330 80 -313
rect 97 -330 105 -313
rect 160 -319 198 -302
rect 72 -338 105 -330
rect 125 -353 158 -345
rect 125 -357 133 -353
rect 108 -370 133 -357
rect 150 -370 158 -353
rect 108 -378 158 -370
rect 108 -435 125 -378
rect 181 -401 198 -319
rect 72 -443 125 -435
rect 72 -460 80 -443
rect 97 -452 125 -443
rect 144 -418 198 -401
rect 215 -389 248 -381
rect 215 -406 223 -389
rect 240 -406 248 -389
rect 215 -414 248 -406
rect 97 -460 105 -452
rect 72 -468 105 -460
rect 144 -485 161 -418
rect 267 -435 284 -285
rect 179 -443 284 -435
rect 179 -460 187 -443
rect 204 -452 284 -443
rect 204 -460 212 -452
rect 179 -468 212 -460
rect 267 -485 284 -452
rect 36 -493 69 -485
rect 36 -527 44 -493
rect 61 -527 69 -493
rect 36 -535 69 -527
rect 90 -493 123 -485
rect 90 -527 98 -493
rect 115 -527 123 -493
rect 90 -535 123 -527
rect 144 -493 177 -485
rect 144 -527 152 -493
rect 169 -527 177 -493
rect 144 -535 177 -527
rect 197 -493 230 -485
rect 197 -527 205 -493
rect 222 -527 230 -493
rect 197 -552 230 -527
rect 251 -493 284 -485
rect 251 -527 259 -493
rect 276 -527 284 -493
rect 251 -535 284 -527
rect 0 -562 327 -552
rect 0 -590 12 -562
rect 0 -600 327 -590
<< viali >>
rect 15 247 32 264
rect 134 257 151 274
rect 50 192 67 209
rect 103 207 120 224
rect 134 157 151 174
rect 255 253 272 270
rect 428 270 445 287
rect 377 242 394 259
rect 480 236 497 253
rect 413 158 430 175
rect 500 167 517 184
rect 621 251 638 268
rect 550 140 567 157
rect 693 140 710 157
rect 98 -277 115 -193
rect 223 -406 240 -389
rect 98 -527 115 -493
<< metal1 >>
rect 145 301 389 315
rect 145 282 159 301
rect 126 274 159 282
rect 374 295 389 301
rect 374 287 453 295
rect 374 281 428 287
rect 7 264 40 272
rect 7 247 15 264
rect 32 247 40 264
rect 126 263 134 274
rect 7 239 40 247
rect 54 257 134 263
rect 151 257 159 274
rect 247 271 280 278
rect 208 270 280 271
rect 54 249 159 257
rect 183 254 255 270
rect 54 216 70 249
rect 183 232 199 254
rect 247 253 255 254
rect 272 253 280 270
rect 420 270 428 281
rect 445 270 453 287
rect 247 245 280 253
rect 369 259 402 267
rect 420 262 453 270
rect 95 224 199 232
rect 42 209 75 216
rect 42 192 50 209
rect 67 192 75 209
rect 95 207 103 224
rect 120 216 199 224
rect 369 242 377 259
rect 394 242 402 259
rect 369 234 402 242
rect 369 223 386 234
rect 120 207 128 216
rect 243 208 386 223
rect 439 211 453 262
rect 613 268 646 276
rect 613 261 621 268
rect 472 253 621 261
rect 472 236 480 253
rect 497 251 621 253
rect 638 251 646 268
rect 497 243 646 251
rect 497 236 505 243
rect 472 228 505 236
rect 95 199 128 207
rect 439 197 492 211
rect 42 150 75 192
rect 478 192 492 197
rect 478 184 525 192
rect 126 176 159 182
rect 405 176 438 183
rect 478 177 500 184
rect 126 175 438 176
rect 126 174 413 175
rect 126 157 134 174
rect 151 162 413 174
rect 151 157 159 162
rect 126 149 159 157
rect 405 158 413 162
rect 430 158 438 175
rect 492 167 500 177
rect 517 167 525 184
rect 492 159 525 167
rect 405 150 438 158
rect 542 157 718 165
rect 542 140 550 157
rect 567 150 693 157
rect 567 140 575 150
rect 542 132 575 140
rect 685 140 693 150
rect 710 140 718 157
rect 685 132 718 140
rect 90 -193 123 -185
rect 90 -277 98 -193
rect 115 -277 123 -193
rect 90 -285 123 -277
rect 109 -388 123 -285
rect 215 -388 248 -381
rect 109 -389 248 -388
rect 109 -403 223 -389
rect 109 -485 123 -403
rect 215 -406 223 -403
rect 240 -406 248 -389
rect 215 -414 248 -406
rect 90 -493 123 -485
rect 90 -527 98 -493
rect 115 -527 123 -493
rect 90 -535 123 -527
<< labels >>
flabel pdiff 87 366 87 366 1 FreeSerif 8 0 0 0 S$
flabel pdiff 141 366 141 366 1 FreeSerif 8 0 0 0 S$
flabel ndiff 141 90 141 90 1 FreeSerif 8 0 0 0 S$
flabel ndiff 87 90 87 90 1 FreeSerif 8 0 0 0 S$
flabel locali 0 432 790 480 0 FreeSerif 80 0 0 0 VDD!
port 15 nsew
flabel locali 0 0 790 48 0 FreeSerif 80 0 0 0 GND!
port 16 nsew
flabel locali 7 239 40 272 0 FreeSerif 80 0 0 0 D
port 0 nsew
flabel locali 42 150 75 183 0 FreeSerif 80 0 0 0 ~CLK
port 1 nsew
flabel pdiff 453 366 453 366 1 FreeSerif 8 0 0 0 S$
flabel pdiff 507 366 507 366 1 FreeSerif 8 0 0 0 S$
flabel ndiff 507 90 507 90 1 FreeSerif 8 0 0 0 S$
flabel ndiff 453 90 453 90 1 FreeSerif 8 0 0 0 S$
flabel locali 405 183 438 216 0 FreeSerif 80 0 0 0 CLK
port 2 nsew
flabel ndiff 628 90 628 90 1 FreeSerif 8 180 0 0 S$
flabel pdiff 628 365 628 365 1 FreeSerif 8 180 0 0 S$
flabel locali 634 185 667 218 0 FreeSerif 80 0 0 0 Q
port 4 nsew
flabel pdiff 667 365 667 365 1 FreeSerif 8 0 0 0 S$
flabel ndiff 667 90 667 90 1 FreeSerif 8 0 0 0 S$
flabel locali 685 182 718 219 0 FreeSerif 80 0 0 0 ~Q
port 3 nsew
flabel pdiff 225 365 225 365 1 FreeSerif 8 180 0 0 S$
flabel ndiff 225 90 225 90 1 FreeSerif 8 180 0 0 S$
flabel ndiff 264 90 264 90 1 FreeSerif 8 0 0 0 S$
flabel pdiff 264 365 264 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 87 -234 87 -234 1 FreeSerif 8 0 0 0 S$
flabel pdiff 141 -234 141 -234 1 FreeSerif 8 0 0 0 S$
flabel ndiff 141 -510 141 -510 1 FreeSerif 8 0 0 0 S$
flabel ndiff 87 -510 87 -510 1 FreeSerif 8 0 0 0 S$
flabel pdiff 194 -235 194 -235 1 FreeSerif 8 180 0 0 S$
flabel ndiff 194 -510 194 -510 1 FreeSerif 8 180 0 0 S$
flabel ndiff 233 -510 233 -510 1 FreeSerif 8 0 0 0 S$
flabel pdiff 233 -235 233 -235 1 FreeSerif 8 0 0 0 S$
<< end >>
