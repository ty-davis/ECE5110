* NGSPICE file created from func_gen_8_connected.ext - technology: sky130A

.subckt memory_8 word0 word1 word2 word3 word4 word5 word6 word7 word8 word9 word10
+ word11 word12 word13 word14 word15 word16 word17 word18 word19 word20 word21 word22
+ word23 word24 word25 word26 word27 word28 word29 word30 word31 word32 word33 word34
+ word35 word36 word37 word38 word39 word40 word41 word42 word43 word44 word45 word46
+ word47 word48 word49 word50 word51 word52 word53 word54 word55 word56 word57 word58
+ word59 word60 word61 word62 word63 word64 word65 word66 word67 word68 word69 word70
+ word71 word72 word73 word74 word75 word76 word77 word78 word79 word80 word81 word82
+ word83 word84 word85 word86 word87 word88 word89 word90 word91 word92 word93 word94
+ word95 word96 word97 word98 word99 word100 word101 word102 word103 word104 word105
+ word106 word107 word108 word109 word110 word111 word112 word113 word114 word115
+ word116 word117 word118 word119 word120 word121 word122 word123 word124 word125
+ word126 word127 word128 word129 word130 word131 word132 word133 word134 word135
+ word136 word137 word138 word139 word140 word141 word142 word143 word144 word145
+ word146 word147 word148 word149 word150 word151 word152 word153 word154 word155
+ word156 word157 word158 word159 word160 word161 word162 word163 word164 word165
+ word166 word167 word168 word169 word170 word171 word172 word173 word174 word175
+ word176 word177 word178 word179 word180 word181 word182 word183 word184 word185
+ word186 word187 word188 word189 word190 word191 word192 word193 word194 word195
+ word196 word197 word198 word199 word200 word201 word202 word203 word204 word205
+ word206 word207 word208 word209 word210 word211 word212 word213 word214 word215
+ word216 word217 word218 word219 word220 word221 word222 word223 word224 word225
+ word226 word227 word228 word229 word230 word231 word232 word233 word234 word235
+ word236 word237 word238 word239 word240 word241 word242 word243 word244 word245
+ word246 word247 word248 word249 word250 word251 word252 word253 word254 word255
+ word256 word257 word258 word259 word260 word261 word262 word263 word264 word265
+ word266 word267 word268 word269 word270 word271 word272 word273 word274 word275
+ word276 word277 word278 word279 word280 word281 word282 word283 word284 word285
+ word286 word287 word288 word289 word290 word291 word292 word293 word294 word295
+ word296 word297 word298 word299 word300 word301 word302 word303 word304 word305
+ word306 word307 word308 word309 word310 word311 word312 word313 word314 word315
+ word316 word317 word318 word319 word320 word321 word322 word323 word324 word325
+ word326 word327 word328 word329 word330 word331 word332 word333 word334 word335
+ word336 word337 word338 word339 word340 word341 word342 word343 word344 word345
+ word346 word347 word348 word349 word350 word351 word352 word353 word354 word355
+ word356 word357 word358 word359 word360 word361 word362 word363 word364 word365
+ word366 word367 word368 word369 word370 word371 word372 word373 word374 word375
+ word376 word377 word378 word379 word380 word381 word382 word383 word384 word385
+ word386 word387 word388 word389 word390 word391 word392 word393 word394 word395
+ word396 word397 word398 word399 word400 word401 word402 word403 word404 word405
+ word406 word407 word408 word409 word410 word411 word412 word413 word414 word415
+ word416 word417 word418 word419 word420 word421 word422 word423 word424 word425
+ word426 word427 word428 word429 word430 word431 word432 word433 word434 word435
+ word436 word437 word438 word439 word440 word441 word442 word443 word444 word445
+ word446 word447 word448 word449 word450 word451 word452 word453 word454 word455
+ word456 word457 word458 word459 word460 word461 word462 word463 word464 word465
+ word466 word467 word468 word469 word470 word471 word472 word473 word474 word475
+ word476 word477 word478 word479 word480 word481 word482 word483 word484 word485
+ word486 word487 word488 word489 word490 word491 word492 word493 word494 word495
+ word496 word497 word498 word499 word500 word501 word502 word503 word504 word505
+ word506 word507 word508 word509 word510 word511 word512 word513 word514 word515
+ word516 word517 word518 word519 word520 word521 word522 word523 word524 word525
+ word526 word527 word528 word529 word530 word531 word532 word533 word534 word535
+ word536 word537 word538 word539 word540 word541 word542 word543 word544 word545
+ word546 word547 word548 word549 word550 word551 word552 word553 word554 word555
+ word556 word557 word558 word559 word560 word561 word562 word563 word564 word565
+ word566 word567 word568 word569 word570 word571 word572 word573 word574 word575
+ word576 word577 word578 word579 word580 word581 word582 word583 word584 word585
+ word586 word587 word588 word589 word590 word591 word592 word593 word594 word595
+ word596 word597 word598 word599 word600 word601 word602 word603 word604 word605
+ word606 word607 word608 word609 word610 word611 word612 word613 word614 word615
+ word616 word617 word618 word619 word620 word621 word622 word623 word624 word625
+ word626 word627 word628 word629 word630 word631 word632 word633 word634 word635
+ word636 word637 word638 word639 word640 word641 word642 word643 word644 word645
+ word646 word647 word648 word649 word650 word651 word652 word653 word654 word655
+ word656 word657 word658 word659 word660 word661 word662 word663 word664 word665
+ word666 word667 word668 word669 word670 word671 word672 word673 word674 word675
+ word676 word677 word678 word679 word680 word681 word682 word683 word684 word685
+ word686 word687 word688 word689 word690 word691 word692 word693 word694 word695
+ word696 word697 word698 word699 word700 word701 word702 word703 word704 word705
+ word706 word707 word708 word709 word710 word711 word712 word713 word714 word715
+ word716 word717 word718 word719 word720 word721 word722 word723 word724 word725
+ word726 word727 word728 word729 word730 word731 word732 word733 word734 word735
+ word736 word737 word738 word739 word740 word741 word742 word743 word744 word745
+ word746 word747 word748 word749 word750 word751 word752 word753 word754 word755
+ word756 word757 word758 word759 word760 word761 word762 word763 word764 word765
+ word766 word767 word768 word769 word770 word771 word772 word773 word774 word775
+ word776 word777 word778 word779 word780 word781 word782 word783 word784 word785
+ word786 word787 word788 word789 word790 word791 word792 word793 word794 word795
+ word796 word797 word798 word799 word800 word801 word802 word803 word804 word805
+ word806 word807 word808 word809 word810 word811 word812 word813 word814 word815
+ word816 word817 word818 word819 word820 word821 word822 word823 word824 word825
+ word826 word827 word828 word829 word830 word831 word832 word833 word834 word835
+ word836 word837 word838 word839 word840 word841 word842 word843 word844 word845
+ word846 word847 word848 word849 word850 word851 word852 word853 word854 word855
+ word856 word857 word858 word859 word860 word861 word862 word863 word864 word865
+ word866 word867 word868 word869 word870 word871 word872 word873 word874 word875
+ word876 word877 word878 word879 word880 word881 word882 word883 word884 word885
+ word886 word887 word888 word889 word890 word891 word892 word893 word894 word895
+ word896 word897 word898 word899 word900 word901 word902 word903 word904 word905
+ word906 word907 word908 word909 word910 word911 word912 word913 word914 word915
+ word916 word917 word918 word919 word920 word921 word922 word923 word924 word925
+ word926 word927 word928 word929 word930 word931 word932 word933 word934 word935
+ word936 word937 word938 word939 word940 word941 word942 word943 word944 word945
+ word946 word947 word948 word949 word950 word951 word952 word953 word954 word955
+ word956 word957 word958 word959 word960 word961 word962 word963 word964 word965
+ word966 word967 word968 word969 word970 word971 word972 word973 word974 word975
+ word976 word977 word978 word979 word980 word981 word982 word983 word984 word985
+ word986 word987 word988 word989 word990 word991 word992 word993 word994 word995
+ word996 word997 word998 word999 word1000 word1001 word1002 word1003 word1004 word1005
+ word1006 word1007 word1008 word1009 word1010 word1011 word1012 word1013 word1014
+ word1015 word1016 word1017 word1018 word1019 word1020 word1021 word1022 word1023
+ Y7 Y6 Y5 Y4 Y3 Y2 Y1 Y0 GND VDD
X0 Y0 word590 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1 GND word1003 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2 Y3 word702 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3 GND word211 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4 Y3 word270 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X5 Y4 word996 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X6 Y4 word838 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X7 GND word207 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X8 GND word215 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X9 GND word365 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X10 Y0 word424 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X11 Y3 word638 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X12 GND word579 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X13 Y7 word924 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X14 GND word865 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X15 GND word143 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X16 GND word867 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X17 Y5 word808 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X18 Y6 word298 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X19 Y6 word628 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X20 GND word137 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X21 Y4 word320 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X22 Y6 word716 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X23 GND word311 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X24 Y0 word470 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X25 GND word625 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X26 Y0 word248 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X27 GND word403 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X28 GND word913 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X29 Y7 word748 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X30 GND word821 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X31 GND word185 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X32 Y7 word224 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X33 GND word361 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X34 GND word511 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X35 Y4 word632 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X36 GND word691 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X37 GND word623 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X38 GND word169 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X39 GND word329 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X40 Y4 word568 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X41 GND word897 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X42 Y6 word862 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X43 GND word385 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X44 Y3 word736 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X45 GND word167 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X46 Y5 word226 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X47 Y2 word894 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X48 Y1 word376 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X49 Y2 word160 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X50 GND word219 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X51 GND word967 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X52 Y6 word908 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X53 GND word841 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X54 GND word151 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X55 Y7 word370 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X56 GND word583 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X57 Y1 word422 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X58 GND word639 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X59 Y7 word700 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X60 Y7 word148 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X61 Y6 word742 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X62 Y3 word718 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X63 Y2 word324 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X64 Y1 word358 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X65 Y1 word688 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X66 Y3 word882 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X67 GND word313 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X68 Y0 word766 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X69 GND word759 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X70 Y7 word682 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X71 Y2 word818 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X72 GND word699 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X73 GND word795 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X74 Y5 word418 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X75 GND word627 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X76 GND word235 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X77 GND word959 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X78 Y1 word900 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X79 Y0 word912 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X80 GND word677 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X81 GND word285 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X82 GND word435 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X83 GND word217 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X84 Y0 word274 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X85 Y6 word590 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X86 GND word935 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X87 GND word905 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X88 Y5 word878 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X89 GND word207 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X90 GND word365 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X91 Y4 word390 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X92 Y0 word540 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X93 GND word381 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X94 Y7 word710 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X95 GND word143 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X96 GND word953 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X97 GND word775 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X98 GND word597 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X99 GND word983 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X100 GND word887 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X101 GND word165 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X102 GND word315 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X103 Y0 word374 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X104 Y3 word588 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X105 Y3 word156 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X106 Y6 word470 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X107 Y7 word874 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X108 Y5 word758 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X109 Y6 word248 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X110 GND word149 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X111 GND word211 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X112 Y4 word270 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X113 GND word479 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X114 Y4 word702 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X115 GND word261 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X116 Y0 word420 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X117 Y4 word638 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X118 GND word987 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X119 Y0 word198 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X120 Y0 word356 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X121 Y4 word536 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X122 Y7 word856 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X123 Y0 word686 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X124 GND word929 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X125 GND word135 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X126 Y7 word174 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X127 GND word461 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X128 GND word707 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X129 Y6 word978 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X130 GND word221 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X131 Y7 word440 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X132 VDD GND Y5 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X133 GND word847 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X134 Y3 word788 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X135 GND word1005 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X136 Y6 word812 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X137 GND word753 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X138 Y0 word668 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X139 GND word335 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X140 Y1 word428 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X141 GND word647 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X142 Y5 word176 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X143 GND word215 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X144 Y1 word326 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X145 Y2 word844 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X146 Y3 word952 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X147 GND word893 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X148 Y2 word780 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X149 GND word169 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X150 GND word383 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X151 Y5 word380 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X152 Y2 word888 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X153 Y2 word376 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X154 Y5 word158 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X155 Y1 word308 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X156 Y5 word488 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X157 Y1 word206 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X158 GND word583 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X159 GND word151 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X160 GND word481 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X161 Y1 word142 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X162 GND word361 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X163 GND word639 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X164 Y1 word472 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X165 GND word691 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X166 Y1 word804 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X167 Y4 word704 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X168 Y2 word688 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X169 GND word185 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X170 GND word673 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X171 GND word845 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X172 GND word235 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X173 GND word385 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X174 Y0 word1020 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X175 GND word167 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X176 Y3 word226 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X177 GND word885 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X178 Y5 word828 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X179 Y0 word798 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X180 GND word219 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X181 GND word891 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X182 GND word791 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X183 Y4 word732 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X184 Y0 word160 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X185 GND word281 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X186 GND word315 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X187 Y6 word374 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X188 GND word433 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X189 Y0 word490 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X190 Y5 word884 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X191 Y3 word272 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X192 GND word719 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X193 GND word217 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X194 Y4 word998 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X195 GND word903 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X196 Y0 word426 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X197 GND word581 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X198 Y4 word896 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X199 GND word149 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X200 GND word265 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X201 Y0 word324 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X202 GND word479 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X203 Y3 word538 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X204 Y7 word926 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X205 GND word765 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X206 Y6 word198 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X207 GND word925 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X208 GND word873 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X209 Y6 word356 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X210 GND word381 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X211 Y4 word156 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X212 GND word699 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X213 Y0 word306 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X214 GND word461 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X215 Y4 word486 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X216 Y3 word418 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X217 GND word879 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X218 GND word363 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X219 Y0 word572 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X220 GND word693 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X221 GND word411 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X222 Y2 word850 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X223 GND word911 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X224 GND word171 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X225 Y7 word390 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X226 Y5 word450 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X227 Y4 word468 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X228 Y0 word618 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X229 GND word797 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X230 GND word659 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X231 Y6 word920 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X232 GND word955 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X233 Y2 word1014 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X234 Y6 word762 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X235 Y5 word228 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X236 Y1 word378 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X237 Y3 word794 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X238 GND word165 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X239 GND word225 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X240 Y1 word276 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X241 Y5 word284 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X242 GND word733 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X243 Y1 word434 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X244 GND word555 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X245 Y5 word614 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X246 Y3 word902 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X247 GND word221 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X248 GND word153 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X249 Y1 word212 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X250 Y7 word372 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X251 GND word431 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X252 GND word899 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X253 GND word211 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X254 Y7 word702 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X255 GND word389 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X256 Y2 word428 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X257 GND word539 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X258 Y2 word996 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X259 GND word267 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X260 Y1 word258 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X261 GND word533 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X262 Y5 word430 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X263 GND word589 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X264 Y1 word580 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X265 GND word701 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X266 Y2 word308 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X267 GND word367 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X268 Y2 word206 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X269 GND word637 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X270 Y2 word694 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X271 Y2 word142 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X272 GND word135 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X273 GND word413 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X274 Y2 word472 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X275 GND word385 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X276 Y1 word736 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X277 GND word185 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X278 GND word219 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X279 GND word907 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X280 Y6 word160 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X281 Y3 word176 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X282 GND word335 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X283 Y0 word970 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X284 GND word943 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X285 Y1 word1002 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X286 GND word835 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X287 GND word605 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X288 Y0 word748 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X289 GND word169 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X290 GND word999 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X291 GND word841 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X292 GND word383 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X293 GND word777 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X294 GND word167 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X295 Y4 word226 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X296 Y3 word158 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X297 Y0 word376 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X298 Y3 word488 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X299 Y7 word876 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X300 GND word433 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X301 GND word151 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X302 Y3 word544 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X303 GND word875 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X304 GND word723 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X305 Y4 word272 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X306 Y6 word306 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X307 GND word331 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X308 Y0 word422 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X309 GND word481 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X310 GND word263 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X311 GND word759 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X312 Y6 word724 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X313 Y0 word358 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X314 Y4 word538 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X315 GND word917 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X316 Y0 word688 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X317 GND word411 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X318 Y4 word594 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X319 Y7 word858 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X320 GND word235 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X321 Y3 word864 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X322 Y7 word756 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X323 GND word313 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X324 Y1 word504 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X325 GND word829 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X326 GND word463 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X327 Y0 word522 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X328 Y6 word618 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X329 GND word859 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X330 Y2 word800 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X331 GND word699 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X332 Y7 word340 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X333 GND word459 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X334 Y4 word418 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X335 GND word747 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X336 GND word217 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X337 GND word905 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X338 Y6 word870 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X339 Y5 word178 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X340 Y1 word328 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X341 GND word175 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X342 Y5 word234 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X343 GND word171 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X344 Y1 word384 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X345 Y1 word162 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X346 Y7 word322 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X347 GND word381 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X348 GND word975 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X349 GND word591 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X350 Y5 word280 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X351 GND word339 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X352 GND word887 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X353 Y7 word156 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X354 Y2 word276 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X355 Y1 word208 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X356 Y7 word644 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X357 GND word153 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X358 Y2 word212 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X359 Y5 word546 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X360 Y1 word696 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X361 GND word363 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X362 GND word935 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X363 GND word693 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X364 Y0 word774 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X365 Y0 word710 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X366 Y5 word904 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X367 Y0 word874 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X368 Y5 word692 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X369 Y3 word450 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X370 Y1 word788 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X371 GND word135 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X372 GND word169 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X373 Y3 word228 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X374 GND word225 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X375 GND word893 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X376 Y4 word852 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X377 GND word793 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X378 GND word221 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X379 Y6 word376 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X380 GND word555 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X381 GND word945 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X382 Y5 word886 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X383 GND word949 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X384 GND word849 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X385 GND word721 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X386 GND word333 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X387 Y0 word428 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X388 GND word727 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X389 GND word151 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X390 Y4 word176 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X391 Y0 word326 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X392 GND word583 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X393 Y7 word928 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X394 Y4 word898 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X395 GND word267 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X396 GND word605 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X397 GND word639 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X398 Y4 word664 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X399 GND word655 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X400 GND word993 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X401 GND word767 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X402 Y6 word358 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X403 GND word383 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X404 Y5 word986 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X405 GND word825 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X406 Y4 word380 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X407 GND word439 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X408 Y4 word158 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X409 Y0 word308 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X410 GND word367 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X411 GND word701 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X412 GND word463 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X413 GND word867 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X414 Y2 word704 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X415 Y0 word206 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X416 Y4 word544 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X417 GND word637 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X418 Y3 word814 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X419 GND word185 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X420 Y0 word694 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X421 Y0 word142 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X422 GND word245 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X423 Y1 word454 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X424 GND word413 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X425 Y0 word472 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X426 GND word627 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X427 Y2 word750 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X428 GND word913 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X429 GND word715 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X430 GND word229 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X431 Y5 word350 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X432 GND word559 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X433 Y6 word922 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X434 Y5 word128 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X435 GND word167 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X436 Y7 word226 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X437 Y2 word504 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X438 Y6 word820 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X439 Y1 word278 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X440 Y5 word286 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X441 Y1 word436 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X442 Y5 word184 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X443 Y1 word334 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X444 Y5 word616 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X445 GND word791 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X446 GND word433 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X447 GND word331 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X448 GND word901 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X449 GND word391 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X450 Y1 word600 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X451 Y2 word328 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X452 Y2 word896 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X453 GND word861 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X454 GND word837 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X455 Y2 word384 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X456 Y2 word162 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X457 GND word591 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X458 GND word373 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X459 GND word489 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X460 GND word937 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X461 GND word703 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X462 Y1 word480 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X463 GND word699 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X464 Y2 word208 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X465 GND word425 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X466 Y7 word418 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X467 Y2 word696 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X468 GND word687 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X469 GND word295 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X470 Y0 word824 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X471 Y3 word400 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X472 GND word459 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X473 GND word797 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X474 GND word221 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X475 Y3 word178 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X476 Y3 word666 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X477 GND word175 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X478 Y3 word234 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X479 Y1 word902 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X480 GND word843 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X481 GND word171 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X482 GND word895 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X483 Y4 word450 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X484 GND word899 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X485 GND word441 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X486 Y4 word228 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X487 Y3 word280 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X488 Y0 word378 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X489 GND word1013 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X490 GND word225 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X491 Y0 word276 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X492 Y4 word284 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X493 Y7 word878 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X494 Y0 word434 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X495 GND word589 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X496 Y7 word934 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X497 GND word153 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X498 Y0 word212 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X499 Y6 word308 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X500 GND word333 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X501 GND word367 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X502 GND word877 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X503 Y6 word206 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X504 GND word483 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X505 Y7 word712 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X506 Y4 word330 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X507 GND word389 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X508 Y6 word142 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X509 Y0 word258 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X510 GND word317 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X511 Y5 word982 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X512 GND word413 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X513 Y6 word472 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X514 Y4 word596 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X515 Y7 word758 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X516 GND word587 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X517 Y6 word890 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X518 Y3 word764 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X519 GND word135 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X520 Y5 word918 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X521 GND word195 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X522 Y5 word254 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X523 Y1 word404 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X524 Y0 word580 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X525 GND word701 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X526 GND word971 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X527 GND word179 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X528 GND word637 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X529 Y2 word966 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X530 GND word931 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X531 Y6 word872 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X532 Y3 word746 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X533 Y7 word176 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X534 Y5 word236 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X535 Y1 word386 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X536 Y7 word664 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X537 Y5 word134 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X538 GND word741 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X539 Y6 word706 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X540 GND word383 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X541 GND word977 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X542 GND word229 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X543 GND word559 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X544 Y1 word652 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X545 Y3 word910 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X546 GND word161 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X547 Y1 word220 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X548 GND word341 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X549 Y7 word380 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X550 GND word439 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X551 Y2 word948 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X552 Y3 word846 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X553 GND word787 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X554 Y7 word158 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X555 Y2 word436 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X556 GND word811 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X557 Y5 word218 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X558 Y5 word548 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X559 Y7 word646 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X560 Y2 word782 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X561 GND word951 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X562 Y3 word892 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X563 GND word541 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X564 Y2 word600 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X565 Y5 word382 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X566 Y1 word532 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X567 GND word835 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X568 GND word375 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X569 Y1 word864 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X570 GND word487 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X571 Y3 word304 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X572 GND word245 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X573 Y2 word582 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X574 GND word423 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X575 Y2 word480 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X576 GND word747 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X577 Y3 word350 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X578 GND word409 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X579 Y5 word740 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X580 GND word687 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X581 GND word171 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X582 GND word981 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X583 Y1 word744 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X584 Y3 word128 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X585 Y3 word286 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X586 Y0 word504 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X587 GND word915 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X588 Y4 word974 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X589 Y0 word858 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X590 Y3 word184 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X591 Y6 word378 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X592 GND word947 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X593 Y1 word1010 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X594 GND word851 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X595 Y0 word756 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X596 Y4 word400 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X597 GND word153 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X598 Y4 word178 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X599 Y6 word212 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X600 Y0 word328 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X601 GND word175 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X602 Y4 word234 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X603 Y4 word666 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X604 Y0 word384 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X605 Y5 word988 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X606 Y7 word884 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X607 Y0 word162 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X608 GND word317 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X609 Y4 word500 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X610 GND word827 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X611 Y3 word432 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X612 Y0 word650 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X613 GND word735 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X614 GND word373 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X615 GND word489 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X616 GND word703 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X617 Y0 word208 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X618 GND word425 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X619 Y6 word580 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X620 GND word925 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X621 Y3 word816 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X622 Y0 word696 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X623 GND word537 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X624 Y5 word868 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X625 Y5 word204 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X626 Y2 word752 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X627 GND word717 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X628 Y0 word530 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X629 Y1 word290 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X630 GND word231 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X631 GND word569 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X632 GND word129 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X633 GND word857 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X634 Y7 word228 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X635 Y5 word288 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X636 GND word881 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X637 Y6 word822 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X638 GND word225 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X639 Y2 word404 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X640 Y5 word186 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X641 Y1 word336 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X642 Y2 word852 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X643 GND word793 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X644 Y3 word962 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X645 Y4 word692 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X646 Y5 word674 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X647 GND word179 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X648 GND word333 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X649 GND word393 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X650 Y5 word452 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X651 Y1 word170 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X652 Y7 word330 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X653 GND word389 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X654 GND word449 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X655 Y2 word898 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X656 GND word863 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X657 Y3 word796 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X658 Y5 word168 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X659 GND word227 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X660 GND word445 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X661 GND word761 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X662 GND word557 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X663 GND word655 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X664 GND word161 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X665 Y2 word220 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X666 GND word493 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X667 Y6 word968 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X668 Y3 word842 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X669 Y7 word430 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X670 Y2 word550 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X671 GND word643 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X672 GND word273 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X673 Y1 word482 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X674 GND word701 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X675 GND word985 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X676 GND word195 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X677 Y3 word254 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X678 Y0 word826 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X679 GND word523 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X680 GND word819 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X681 Y4 word760 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X682 GND word245 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X683 Y4 word304 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X684 Y0 word454 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X685 Y3 word236 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X686 GND word609 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X687 Y7 word954 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X688 Y3 word134 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X689 GND word573 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X690 Y0 word808 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X691 GND word901 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X692 GND word897 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X693 Y4 word860 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X694 GND word229 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X695 GND word443 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X696 Y5 word894 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X697 Y4 word350 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X698 Y6 word384 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X699 GND word729 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X700 Y4 word128 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X701 Y6 word162 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X702 GND word341 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X703 GND word499 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X704 Y0 word278 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X705 Y4 word286 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X706 Y0 word436 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X707 GND word495 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X708 Y4 word184 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X709 Y3 word218 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X710 Y0 word334 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X711 GND word591 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X712 Y7 word936 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X713 GND word965 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X714 Y4 word906 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X715 GND word607 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X716 Y1 word942 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X717 Y7 word834 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X718 VDD GND Y7 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X719 Y6 word208 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X720 GND word391 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X721 Y5 word994 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X722 Y3 word382 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X723 Y0 word600 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X724 GND word711 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X725 Y4 word598 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X726 GND word657 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X727 Y1 word140 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X728 GND word375 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X729 GND word875 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X730 Y3 word766 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X731 Y7 word354 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X732 Y4 word432 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X733 Y0 word582 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X734 Y6 word726 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X735 GND word703 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X736 Y0 word480 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X737 GND word181 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X738 Y1 word240 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X739 Y7 word400 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X740 GND word537 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X741 GND word933 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X742 Y7 word178 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X743 Y3 word866 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X744 Y5 word238 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X745 GND word831 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X746 Y5 word136 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X747 GND word175 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X748 Y7 word234 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X749 Y7 word666 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X750 GND word743 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X751 Y6 word708 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X752 GND word231 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X753 Y5 word624 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X754 GND word129 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X755 Y1 word222 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X756 GND word441 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X757 GND word339 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X758 GND word343 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X759 Y1 word552 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X760 GND word399 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X761 GND word497 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X762 Y2 word1006 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X763 GND word813 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X764 GND word177 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X765 Y2 word336 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X766 Y2 word170 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X767 Y1 word368 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X768 GND word275 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X769 Y1 word764 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X770 Y3 word204 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X771 Y0 word878 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X772 Y6 word454 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X773 Y0 word934 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X774 Y5 word964 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X775 Y7 word692 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X776 GND word569 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X777 Y0 word712 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X778 GND word983 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X779 GND word195 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X780 GND word229 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X781 Y4 word254 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X782 Y3 word288 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X783 Y0 word404 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X784 GND word739 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X785 Y3 word186 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X786 Y7 word904 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X787 Y0 word758 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X788 Y4 word810 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X789 GND word179 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X790 GND word393 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X791 Y5 word844 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X792 Y1 word846 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X793 GND word787 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X794 GND word449 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X795 Y4 word236 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X796 Y0 word386 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X797 GND word445 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X798 Y6 word600 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X799 Y4 word134 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X800 Y3 word168 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X801 GND word227 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X802 GND word945 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X803 Y7 word886 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X804 GND word557 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X805 Y5 word888 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X806 Y4 word502 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X807 Y0 word652 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X808 GND word951 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X809 Y1 word892 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X810 Y4 word792 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X811 GND word161 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X812 Y0 word220 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X813 GND word375 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X814 Y0 word550 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X815 Y5 word944 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X816 GND word491 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X817 GND word499 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X818 Y7 word720 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X819 Y4 word218 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X820 GND word427 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X821 Y6 word582 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X822 GND word607 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X823 GND word325 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X824 GND word927 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X825 GND word245 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X826 Y4 word382 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X827 Y0 word532 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X828 GND word869 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X829 Y2 word140 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X830 GND word131 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X831 Y1 word190 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X832 Y7 word350 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X833 GND word409 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X834 GND word487 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X835 GND word619 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X836 GND word883 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X837 Y7 word128 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X838 Y2 word974 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X839 Y5 word188 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X840 GND word247 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X841 Y6 word880 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X842 Y7 word184 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X843 GND word423 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X844 Y5 word244 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X845 Y1 word394 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X846 GND word181 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X847 Y2 word240 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X848 GND word749 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X849 Y1 word172 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X850 GND word391 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X851 Y1 word660 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X852 GND word349 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X853 Y2 word956 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X854 GND word763 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X855 Y1 word438 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X856 GND word657 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X857 Y1 word494 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X858 Y5 word556 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X859 GND word615 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X860 Y2 word222 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X861 GND word903 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X862 GND word213 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X863 GND word373 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X864 Y7 word432 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X865 Y2 word552 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X866 Y0 word1004 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X867 GND word543 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X868 GND word549 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X869 GND word703 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X870 GND word599 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X871 GND word327 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X872 Y1 word318 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X873 Y1 word816 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X874 GND word779 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X875 GND word809 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X876 Y0 word828 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X877 GND word821 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X878 Y6 word404 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X879 Y5 word914 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X880 Y2 word368 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X881 Y5 word850 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X882 GND word755 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X883 GND word179 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X884 Y4 word204 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X885 Y3 word238 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X886 Y3 word136 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X887 Y3 word294 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X888 GND word473 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X889 Y3 word624 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X890 Y4 word862 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X891 GND word231 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X892 Y0 word290 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X893 Y6 word386 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X894 GND word569 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X895 GND word129 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X896 GND word343 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X897 Y3 word402 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X898 GND word731 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X899 Y4 word288 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X900 GND word497 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X901 Y4 word908 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X902 GND word161 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X903 Y4 word186 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X904 Y6 word220 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X905 Y0 word336 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X906 GND word395 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X907 GND word177 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X908 GND word895 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X909 Y7 word836 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X910 GND word665 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X911 Y4 word452 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X912 Y0 word602 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X913 Y1 word842 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X914 Y0 word170 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X915 GND word449 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X916 GND word227 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X917 Y4 word168 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X918 GND word377 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X919 GND word275 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X920 GND word985 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X921 GND word877 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X922 VDD GND Y2 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X923 GND word195 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X924 Y7 word254 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X925 Y5 word314 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X926 Y4 word332 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X927 Y1 word464 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X928 Y0 word482 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X929 Y6 word728 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X930 Y2 word760 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X931 GND word725 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X932 GND word239 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X933 GND word419 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X934 Y7 word918 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X935 VDD GND Y3 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X936 GND word865 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X937 Y5 word138 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X938 GND word197 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X939 Y7 word236 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X940 GND word889 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X941 Y6 word830 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X942 Y7 word134 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X943 Y1 word564 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X944 Y5 word626 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X945 GND word685 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X946 Y5 word194 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X947 Y1 word344 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X948 GND word131 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X949 Y2 word190 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X950 GND word443 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X951 GND word341 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X952 Y5 word460 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X953 Y3 word748 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X954 Y7 word218 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X955 GND word397 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X956 Y6 word930 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X957 Y1 word388 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X958 Y1 word444 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X959 Y2 word172 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X960 GND word163 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X961 GND word323 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X962 Y7 word382 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X963 GND word651 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X964 Y7 word648 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X965 Y1 word268 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X966 GND word759 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X967 GND word213 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X968 GND word423 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X969 GND word543 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X970 GND word995 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X971 GND word599 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X972 GND word929 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X973 Y0 word140 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X974 Y1 word866 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X975 GND word807 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X976 Y6 word290 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X977 Y5 word800 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X978 GND word231 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X979 GND word247 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X980 GND word129 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X981 Y3 word188 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X982 Y3 word244 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X983 Y0 word240 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X984 GND word753 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X985 GND word181 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X986 GND word395 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X987 GND word905 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X988 Y7 word740 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X989 Y4 word238 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X990 GND word297 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X991 GND word349 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X992 GND word447 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X993 Y6 word602 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X994 Y4 word136 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X995 Y6 word170 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X996 GND word345 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X997 GND word947 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X998 Y0 word980 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X999 GND word853 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1000 Y0 word222 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1001 Y3 word556 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1002 Y5 word946 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1003 GND word887 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1004 GND word377 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1005 Y4 word402 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1006 Y0 word552 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1007 Y7 word722 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1008 Y6 word854 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1009 GND word159 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1010 GND word177 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1011 GND word327 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1012 GND word665 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1013 Y3 word656 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1014 GND word935 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1015 GND word987 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1016 Y6 word900 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1017 Y7 word204 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1018 Y1 word414 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1019 Y6 word734 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1020 GND word133 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1021 Y0 word368 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1022 Y7 word868 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1023 Y0 word698 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1024 GND word189 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1025 Y2 word976 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1026 Y7 word186 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1027 Y2 word464 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1028 Y3 word874 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1029 GND word815 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1030 Y5 word246 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1031 GND word305 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1032 GND word473 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1033 Y7 word674 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1034 Y2 word810 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1035 GND word751 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1036 GND word233 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1037 GND word239 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1038 GND word393 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1039 GND word571 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1040 Y1 word230 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1041 GND word351 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1042 Y1 word560 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1043 Y7 word168 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1044 GND word227 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1045 GND word347 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1046 GND word505 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1047 GND word287 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1048 Y1 word338 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1049 Y1 word496 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1050 GND word283 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1051 Y2 word344 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1052 GND word617 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1053 Y2 word792 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1054 Y5 word676 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1055 GND word961 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X1056 GND word669 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1057 Y7 word332 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1058 Y5 word392 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1059 GND word451 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1060 Y0 word904 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X1061 Y2 word388 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1062 Y2 word444 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1063 Y6 word140 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1064 GND word163 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1065 Y5 word704 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1066 GND word945 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X1067 Y0 word886 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1068 GND word879 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1069 Y2 word268 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1070 GND word419 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1071 GND word181 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1072 Y6 word240 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1073 Y5 word750 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1074 Y0 word720 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1075 GND word197 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1076 Y4 word364 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1077 Y3 word138 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1078 Y4 word984 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1079 GND word685 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1080 Y3 word194 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1081 GND word131 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1082 Y0 word190 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1083 Y4 word762 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1084 GND word469 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1085 GND word401 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1086 Y4 word188 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1087 Y6 word222 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1088 GND word247 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1089 GND word397 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1090 Y4 word244 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1091 Y0 word394 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1092 GND word897 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1093 GND word667 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1094 Y7 word894 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1095 Y1 word154 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1096 Y0 word172 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1097 Y5 word896 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1098 Y0 word660 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1099 GND word349 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1100 Y3 word442 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1101 GND word745 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1102 Y0 word438 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1103 GND word593 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1104 Y7 word938 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1105 GND word277 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1106 Y0 word494 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1107 GND word885 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1108 Y3 word606 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1109 GND word909 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1110 GND word213 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1111 Y5 word316 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1112 Y6 word368 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1113 GND word821 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X1114 GND word713 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1115 GND word719 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1116 Y5 word150 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1117 Y1 word300 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1118 Y0 word318 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1119 GND word421 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1120 GND word139 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1121 GND word473 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1122 Y3 word926 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1123 Y7 word238 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1124 GND word891 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1125 Y7 word136 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1126 GND word765 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1127 Y5 word196 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1128 GND word255 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1129 Y2 word862 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1130 GND word133 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1131 GND word183 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1132 Y7 word402 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1133 GND word189 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1134 GND word343 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1135 Y5 word462 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1136 Y1 word180 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1137 GND word399 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1138 Y1 word612 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1139 GND word671 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1140 Y6 word932 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1141 GND word873 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1142 GND word177 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1143 GND word237 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1144 Y1 word446 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1145 GND word665 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1146 GND word233 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1147 Y2 word742 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1148 Y2 word230 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1149 Y5 word342 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1150 Y2 word560 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1151 GND word159 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1152 Y1 word492 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1153 GND word551 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1154 Y2 word496 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1155 Y4 word724 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1156 Y3 word264 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1157 Y2 word542 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1158 GND word997 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1159 Y1 word592 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1160 GND word895 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1161 GND word829 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1162 Y1 word924 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X1163 Y5 word802 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1164 GND word131 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1165 Y6 word190 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1166 Y4 word314 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1167 Y0 word464 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1168 GND word619 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1169 Y3 word246 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1170 GND word397 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1171 Y5 word966 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1172 GND word907 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1173 GND word877 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1174 GND word239 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1175 Y6 word394 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1176 GND word419 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1177 GND word571 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1178 GND word351 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1179 Y3 word410 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1180 Y1 word748 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1181 GND word739 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1182 Y4 word138 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1183 Y6 word172 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1184 GND word197 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1185 GND word347 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1186 GND word741 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1187 GND word505 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1188 Y0 word564 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1189 Y4 word626 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1190 GND word975 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1191 Y4 word194 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1192 GND word287 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1193 Y0 word344 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1194 GND word617 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1195 Y0 word918 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X1196 GND word283 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1197 Y5 word948 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1198 GND word1011 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X1199 Y7 word844 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1200 GND word401 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1201 Y0 word610 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1202 Y3 word392 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1203 GND word451 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1204 Y6 word754 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1205 GND word213 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1206 Y0 word388 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1207 GND word209 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1208 Y7 word888 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1209 GND word667 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1210 Y2 word154 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1211 Y0 word444 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1212 GND word599 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1213 GND word835 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1214 Y7 word944 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1215 GND word145 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1216 GND word163 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1217 Y6 word318 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1218 Y7 word364 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1219 GND word501 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1220 GND word929 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1221 Y6 word736 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1222 GND word259 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1223 Y1 word250 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1224 Y0 word268 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1225 Y4 word606 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1226 Y7 word188 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1227 GND word247 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1228 GND word307 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1229 Y1 word516 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1230 GND word205 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1231 Y7 word244 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1232 GND word359 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1233 Y6 word718 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1234 GND word141 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1235 Y2 word300 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1236 GND word139 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1237 Y1 word232 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1238 Y5 word570 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1239 Y1 word130 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1240 GND word349 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1241 GND word917 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X1242 Y3 word858 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1243 Y2 word566 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1244 Y6 word882 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1245 GND word823 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1246 GND word405 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1247 Y1 word498 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1248 Y5 word678 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1249 GND word187 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1250 Y1 word396 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1251 GND word853 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1252 GND word183 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1253 GND word675 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1254 GND word671 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1255 Y2 word180 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1256 GND word453 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1257 GND word603 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1258 Y2 word958 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X1259 GND word923 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1260 Y0 word740 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1261 Y5 word558 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1262 Y7 word656 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1263 GND word653 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1264 Y2 word492 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1265 GND word551 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1266 GND word947 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1267 GND word159 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1268 GND word309 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1269 Y4 word940 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1270 Y3 word150 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1271 Y6 word464 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1272 Y0 word722 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1273 Y5 word752 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1274 GND word357 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1275 GND word239 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1276 Y0 word414 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1277 Y0 word988 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1278 Y3 word196 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1279 GND word255 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1280 Y2 word592 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1281 Y7 word914 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1282 GND word133 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1283 GND word979 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1284 GND word471 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1285 Y7 word850 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1286 Y4 word820 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1287 GND word189 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1288 GND word521 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1289 Y5 word852 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1290 Y1 word856 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1291 Y4 word246 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1292 Y0 word514 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1293 GND word849 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1294 GND word237 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1295 Y3 word296 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1296 GND word455 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1297 Y6 word610 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1298 GND word955 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1299 GND word233 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1300 Y6 word388 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1301 GND word571 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1302 Y5 word898 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1303 GND word861 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1304 Y0 word230 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1305 GND word289 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1306 GND word733 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1307 GND word351 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1308 Y0 word560 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1309 Y7 word730 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1310 Y3 word342 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1311 GND word163 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1312 GND word287 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1313 Y0 word338 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1314 Y0 word496 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1315 Y7 word838 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1316 Y3 word608 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1317 GND word451 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1318 Y0 word542 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1319 Y5 word152 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1320 GND word879 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1321 GND word209 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1322 Y1 word302 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1323 Y5 word640 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1324 Y1 word200 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1325 GND word419 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1326 Y3 word928 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1327 Y4 word658 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1328 GND word145 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1329 GND word893 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1330 Y3 word826 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1331 GND word767 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1332 Y7 word138 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1333 GND word197 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1334 GND word355 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1335 Y1 word466 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1336 GND word685 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1337 Y7 word194 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1338 Y0 word642 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1339 GND word727 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1340 Y2 word250 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1341 Y1 word182 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1342 GND word241 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1343 GND word401 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1344 Y3 word808 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1345 GND word457 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1346 Y1 word448 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1347 Y5 word628 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1348 GND word667 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1349 GND word137 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1350 Y1 word346 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1351 GND word803 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1352 Y2 word232 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1353 GND word291 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1354 GND word625 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1355 Y3 word972 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1356 Y5 word684 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1357 GND word223 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1358 Y1 word282 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1359 Y7 word442 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1360 GND word621 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1361 Y2 word130 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1362 Y2 word396 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1363 GND word885 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1364 Y0 word154 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1365 GND word309 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1366 GND word897 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1367 GND word719 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1368 Y2 word662 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1369 Y4 word890 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1370 GND word259 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1371 Y0 word894 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1372 Y6 word414 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1373 GND word437 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1374 GND word759 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1375 Y1 word926 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X1376 GND word133 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1377 Y4 word316 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1378 GND word919 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1379 Y1 word824 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1380 GND word189 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1381 Y3 word366 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1382 GND word205 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1383 Y0 word938 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1384 GND word931 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1385 Y4 word150 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1386 Y0 word300 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1387 GND word359 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1388 Y0 word994 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1389 GND word139 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1390 GND word141 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1391 GND word421 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1392 GND word455 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1393 GND word859 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1394 GND word233 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1395 Y3 word570 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1396 GND word743 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1397 Y0 word566 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1398 Y4 word196 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1399 Y6 word230 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1400 GND word255 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1401 GND word289 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1402 GND word799 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1403 GND word187 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1404 GND word405 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1405 GND word183 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1406 GND word905 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1407 Y0 word818 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X1408 GND word911 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X1409 Y0 word180 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1410 Y0 word612 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1411 GND word159 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1412 GND word237 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1413 GND word387 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1414 Y0 word446 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1415 GND word601 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1416 Y7 word946 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1417 GND word887 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1418 GND word147 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1419 Y3 word558 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1420 GND word503 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1421 Y6 word738 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1422 Y0 word492 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1423 GND word829 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X1424 Y1 word252 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1425 Y4 word608 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1426 Y3 word934 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1427 Y6 word902 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1428 GND word207 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1429 Y7 word246 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1430 GND word899 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1431 Y1 word416 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1432 Y5 word424 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1433 Y0 word592 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1434 GND word983 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1435 Y2 word870 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1436 GND word695 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1437 GND word143 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1438 Y2 word200 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1439 Y1 word352 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1440 GND word191 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1441 Y7 word410 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1442 Y1 word132 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1443 GND word351 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1444 GND word679 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1445 Y5 word248 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1446 Y1 word398 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1447 Y7 word676 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1448 Y2 word182 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1449 GND word241 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1450 GND word173 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1451 Y7 word392 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1452 Y6 word154 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1453 Y0 word964 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1454 Y2 word448 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1455 Y7 word658 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1456 GND word735 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1457 GND word223 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1458 Y4 word840 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1459 Y3 word152 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1460 GND word209 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1461 Y0 word844 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X1462 Y3 word640 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1463 GND word783 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X1464 Y0 word780 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1465 GND word145 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1466 Y4 word266 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1467 Y6 word300 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1468 GND word359 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1469 GND word869 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1470 Y7 word704 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1471 GND word139 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1472 Y0 word888 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1473 GND word881 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1474 Y0 word250 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1475 GND word405 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1476 GND word915 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1477 GND word917 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X1478 Y1 word858 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1479 Y7 word750 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1480 GND word183 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1481 GND word851 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1482 Y4 word366 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1483 GND word457 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1484 Y0 word516 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1485 Y1 word756 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1486 Y6 word180 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1487 GND word205 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1488 Y6 word612 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1489 GND word957 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1490 GND word749 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1491 GND word137 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1492 GND word141 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1493 GND word963 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1494 GND word863 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1495 Y3 word684 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1496 Y0 word232 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1497 GND word291 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1498 GND word387 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1499 GND word761 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1500 Y0 word130 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1501 GND word403 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1502 Y0 word562 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1503 Y4 word570 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1504 Y7 word732 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1505 Y6 word864 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1506 Y0 word498 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1507 GND word187 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1508 GND word337 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1509 Y0 word396 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1510 Y3 word1004 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1511 Y7 word896 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1512 GND word837 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1513 GND word969 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1514 GND word453 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1515 Y0 word662 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1516 Y5 word274 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1517 Y2 word940 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1518 GND word747 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1519 Y7 word150 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1520 Y1 word202 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1521 GND word421 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1522 Y6 word744 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1523 GND word437 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1524 Y6 word592 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1525 GND word147 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1526 GND word937 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1527 GND word357 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1528 Y3 word884 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1529 Y7 word196 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1530 GND word255 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1531 GND word315 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1532 Y5 word374 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1533 Y1 word524 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1534 Y2 word922 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1535 Y2 word252 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1536 GND word243 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1537 GND word149 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1538 Y5 word420 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1539 Y2 word416 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1540 Y5 word198 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1541 GND word237 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1542 Y2 word574 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1543 GND word809 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X1544 Y1 word348 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1545 Y1 word506 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1546 Y5 word686 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1547 Y2 word352 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1548 Y2 word132 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1549 GND word191 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1550 Y7 word342 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1551 GND word679 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1552 GND word461 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1553 GND word611 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1554 Y0 word914 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1555 GND word209 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1556 GND word173 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1557 GND word145 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1558 GND word661 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1559 GND word955 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X1560 GND word985 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1561 Y1 word928 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X1562 Y3 word590 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1563 GND word921 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1564 GND word789 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X1565 GND word767 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X1566 Y0 word730 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1567 Y4 word726 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1568 Y6 word250 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1569 Y5 word760 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1570 GND word207 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1571 GND word365 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1572 Y3 word424 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1573 Y4 word152 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1574 Y0 word996 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1575 GND word143 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1576 Y0 word302 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1577 GND word457 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1578 Y4 word640 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1579 GND word831 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1580 Y0 word200 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1581 GND word801 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1582 Y6 word232 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1583 GND word291 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1584 GND word407 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1585 Y0 word466 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1586 GND word621 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1587 Y6 word130 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1588 Y3 word248 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1589 GND word907 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1590 GND word709 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1591 Y1 word972 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X1592 Y0 word182 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1593 GND word241 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1594 Y6 word396 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1595 GND word965 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1596 Y5 word906 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1597 GND word741 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1598 Y4 word298 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1599 Y6 word814 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1600 Y0 word448 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1601 GND word507 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1602 GND word603 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1603 Y4 word628 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1604 GND word137 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1605 Y0 word346 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1606 Y7 word948 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1607 GND word625 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1608 Y0 word282 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1609 GND word223 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1610 GND word385 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1611 GND word403 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1612 Y2 word890 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1613 GND word855 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1614 GND word723 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1615 GND word729 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1616 Y5 word160 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1617 GND word219 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1618 Y5 word490 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1619 Y7 word366 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1620 GND word995 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X1621 Y5 word426 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1622 GND word901 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1623 Y1 word144 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1624 GND word205 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1625 Y1 word576 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1626 GND word635 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1627 Y1 word474 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1628 GND word141 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1629 Y2 word202 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1630 GND word193 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1631 Y7 word412 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1632 GND word249 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1633 GND word977 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1634 GND word875 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1635 Y7 word678 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1636 GND word187 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1637 Y5 word306 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1638 Y1 word456 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1639 GND word515 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1640 GND word675 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1641 GND word243 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1642 GND word299 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1643 Y5 word572 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1644 GND word629 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1645 Y1 word620 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1646 Y2 word348 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1647 GND word565 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1648 Y0 word800 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X1649 Y5 word618 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1650 GND word677 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1651 GND word435 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1652 Y2 word670 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1653 Y1 word878 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1654 GND word147 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1655 Y3 word540 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1656 GND word871 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1657 Y6 word302 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1658 Y1 word934 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1659 Y6 word200 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1660 Y3 word374 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1661 Y1 word712 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1662 GND word983 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X1663 GND word883 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1664 Y0 word252 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1665 GND word407 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1666 Y6 word466 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1667 GND word939 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X1668 Y4 word880 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1669 Y7 word752 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1670 GND word149 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1671 GND word817 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X1672 Y5 word810 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1673 GND word751 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1674 Y6 word182 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1675 GND word207 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1676 GND word241 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1677 GND word365 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1678 Y0 word416 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1679 Y0 word574 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1680 Y3 word198 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1681 GND word695 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1682 GND word143 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1683 GND word293 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1684 Y0 word352 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1685 GND word987 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1686 Y3 word686 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1687 GND word191 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1688 Y6 word448 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1689 Y7 word852 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1690 GND word763 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1691 Y0 word132 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1692 Y4 word470 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1693 GND word529 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1694 GND word849 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1695 Y6 word764 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1696 GND word223 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1697 Y4 word248 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1698 Y0 word398 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1699 GND word735 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1700 Y7 word898 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1701 GND word971 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1702 Y3 word904 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1703 Y3 word668 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1704 GND word173 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1705 Y1 word214 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1706 VDD GND Y0 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X1707 Y7 word152 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1708 Y6 word746 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1709 GND word169 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1710 GND word717 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1711 Y1 word260 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1712 GND word945 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X1713 Y3 word886 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1714 Y5 word376 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1715 Y6 word910 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1716 GND word881 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1717 Y3 word720 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1718 GND word151 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1719 Y1 word360 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1720 GND word199 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1721 Y5 word422 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1722 GND word481 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1723 GND word631 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1724 GND word639 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1725 GND word927 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1726 Y2 word576 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1727 Y6 word892 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1728 Y2 word144 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1729 GND word567 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1730 GND word825 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1731 GND word137 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1732 GND word863 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1733 Y5 word688 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1734 Y1 word406 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1735 Y7 word684 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1736 GND word193 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1737 Y0 word704 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1738 GND word249 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1739 GND word403 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1740 GND word463 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1741 Y1 word672 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1742 Y2 word968 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1743 Y2 word456 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1744 Y1 word1004 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1745 Y0 word750 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1746 GND word627 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1747 GND word385 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1748 GND word147 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1749 GND word957 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X1750 Y4 word950 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1751 Y3 word160 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1752 GND word219 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1753 Y3 word490 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1754 Y1 word828 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1755 Y4 word728 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1756 Y6 word252 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1757 Y0 word732 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1758 GND word435 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1759 Y1 word884 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1760 GND word725 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1761 Y3 word426 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1762 Y0 word998 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1763 Y0 word202 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1764 Y0 word896 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1765 GND word837 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X1766 Y4 word540 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1767 GND word889 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1768 Y4 word830 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1769 GND word919 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1770 GND word293 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1771 GND word191 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1772 Y6 word132 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1773 GND word315 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1774 Y0 word524 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1775 GND word243 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1776 GND word967 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1777 Y5 word908 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1778 GND word149 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1779 Y6 word398 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1780 Y4 word930 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1781 GND word743 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1782 GND word299 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1783 Y4 word420 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1784 Y3 word572 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1785 Y6 word816 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1786 GND word411 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1787 GND word173 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1788 Y4 word198 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1789 Y5 word742 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1790 Y0 word348 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1791 Y0 word506 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1792 Y3 word618 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1793 Y1 word164 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1794 Y6 word916 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1795 GND word857 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1796 GND word731 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1797 Y0 word670 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1798 GND word755 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1799 GND word221 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1800 Y1 word210 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1801 GND word997 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1802 Y2 word726 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1803 Y4 word668 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1804 Y6 word962 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1805 GND word895 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1806 GND word207 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1807 Y2 word214 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1808 Y5 word428 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1809 GND word485 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1810 Y3 word836 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1811 Y1 word146 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1812 GND word365 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1813 Y7 word424 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1814 Y1 word476 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1815 GND word535 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1816 GND word933 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X1817 GND word695 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1818 GND word831 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X1819 GND word143 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1820 GND word989 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1821 GND word737 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1822 Y2 word260 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1823 GND word319 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1824 GND word251 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1825 Y1 word310 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1826 Y7 word248 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1827 Y2 word526 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1828 Y5 word308 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1829 Y5 word206 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1830 GND word813 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X1831 GND word697 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1832 Y5 word694 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1833 Y5 word142 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1834 Y2 word360 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1835 Y3 word982 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1836 GND word199 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1837 Y1 word292 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1838 GND word631 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1839 GND word563 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1840 Y3 word918 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1841 GND word567 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1842 GND word465 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1843 Y1 word954 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X1844 GND word795 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1845 GND word335 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1846 Y2 word672 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1847 Y0 word966 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1848 GND word663 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1849 Y4 word900 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1850 GND word169 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1851 Y1 word936 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X1852 GND word995 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X1853 Y6 word202 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1854 Y1 word834 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1855 GND word385 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1856 Y4 word734 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1857 Y3 word376 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1858 Y0 word948 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1859 GND word1007 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X1860 GND word711 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1861 Y4 word160 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1862 GND word219 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1863 GND word941 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1864 Y4 word1000 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1865 GND word151 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1866 GND word369 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1867 GND word839 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1868 GND word481 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1869 GND word639 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1870 GND word869 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1871 Y0 word782 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1872 GND word243 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1873 GND word875 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X1874 GND word753 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1875 Y0 word144 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1876 Y0 word576 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1877 GND word265 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1878 GND word299 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1879 Y3 word358 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1880 GND word415 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1881 Y0 word474 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1882 GND word629 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1883 Y3 word688 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1884 GND word915 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1885 GND word193 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1886 GND word531 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1887 Y1 word980 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1888 GND word851 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1889 GND word249 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1890 Y3 word522 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1891 GND word853 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1892 Y6 word766 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1893 GND word749 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1894 Y0 word456 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1895 GND word611 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1896 Y7 word956 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1897 Y1 word216 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1898 GND word435 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1899 Y4 word572 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1900 Y0 word620 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1901 Y6 word866 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1902 GND word171 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1903 Y2 word778 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1904 VDD GND Y1 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X1905 Y2 word164 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1906 Y6 word912 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1907 GND word155 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1908 Y7 word374 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1909 Y5 word378 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1910 Y5 word276 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1911 Y1 word584 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1912 GND word153 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1913 Y5 word212 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1914 GND word371 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1915 GND word939 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X1916 Y2 word880 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1917 GND word149 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1918 Y2 word210 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1919 Y1 word362 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1920 GND word483 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1921 GND word201 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1922 Y7 word420 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1923 Y3 word988 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1924 Y2 word146 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1925 Y7 word198 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1926 Y7 word356 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1927 Y2 word476 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X1928 GND word535 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1929 GND word317 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1930 Y1 word408 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1931 Y7 word686 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1932 GND word251 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1933 Y1 word242 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1934 GND word517 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X1935 Y0 word752 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1936 Y1 word508 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X1937 Y7 word668 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1938 Y2 word292 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X1939 GND word973 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X1940 Y2 word622 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1941 GND word781 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1942 GND word221 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1943 GND word909 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1944 GND word793 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1945 Y1 word886 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1946 Y0 word214 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1947 GND word335 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1948 GND word369 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1949 GND word879 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1950 GND word849 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X1951 GND word485 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1952 Y7 word714 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1953 Y3 word326 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X1954 GND word663 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1955 Y0 word898 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1956 Y1 word720 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X1957 Y6 word144 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1958 GND word169 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1959 GND word319 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1960 GND word635 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1961 GND word921 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1962 GND word891 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1963 Y0 word260 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1964 GND word415 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X1965 Y6 word474 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1966 Y5 word984 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1967 GND word589 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1968 Y7 word760 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1969 GND word193 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1970 Y5 word920 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1971 GND word825 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X1972 Y5 word762 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1973 GND word367 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X1974 Y0 word526 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1975 GND word249 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1976 GND word697 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X1977 Y3 word206 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1978 Y4 word932 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X1979 GND word151 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1980 GND word301 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1981 Y0 word360 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1982 Y3 word142 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1983 Y4 word422 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1984 Y6 word456 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1985 GND word481 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1986 GND word639 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1987 Y7 word860 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1988 Y0 word690 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X1989 GND word199 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1990 Y3 word472 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X1991 GND word803 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X1992 Y0 word406 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X1993 GND word465 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X1994 Y6 word620 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X1995 Y1 word166 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1996 GND word385 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X1997 Y7 word906 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X1998 Y0 word672 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X1999 Y2 word950 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2000 GND word757 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2001 Y7 word160 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2002 GND word219 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2003 GND word609 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2004 Y2 word728 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2005 Y2 word216 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2006 GND word627 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2007 GND word897 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2008 GND word725 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2009 Y7 word426 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2010 Y7 word324 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2011 Y1 word478 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2012 Y3 word894 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2013 Y5 word384 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2014 Y5 word162 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2015 GND word889 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2016 GND word253 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2017 Y1 word312 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2018 GND word155 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2019 GND word489 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2020 GND word903 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2021 Y2 word584 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2022 Y5 word208 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2023 GND word425 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2024 GND word575 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2025 GND word713 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2026 Y2 word930 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X2027 Y5 word696 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2028 GND word201 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2029 GND word683 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2030 Y1 word192 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2031 GND word411 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2032 Y1 word680 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2033 Y2 word408 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2034 Y1 word458 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2035 GND word919 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2036 Y4 word754 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2037 GND word677 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2038 Y2 word242 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2039 Y1 word790 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X2040 GND word731 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2041 Y6 word214 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2042 GND word171 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2043 Y2 word508 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X2044 GND word997 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2045 Y5 word990 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2046 GND word895 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2047 Y4 word736 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2048 Y0 word164 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2049 GND word319 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2050 GND word829 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2051 GND word799 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2052 Y3 word434 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2053 GND word613 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2054 GND word943 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2055 Y4 word1002 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2056 GND word221 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2057 GND word371 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2058 GND word585 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2059 GND word153 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2060 Y0 word210 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2061 Y3 word212 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2062 GND word269 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2063 GND word999 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2064 GND word871 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2065 GND word841 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2066 GND word483 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2067 GND word539 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2068 Y0 word146 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2069 GND word267 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2070 GND word301 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2071 Y6 word360 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2072 Y5 word870 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2073 GND word199 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2074 GND word317 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2075 Y0 word476 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2076 GND word631 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2077 GND word705 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2078 GND word533 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2079 Y1 word982 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X2080 Y4 word882 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2081 GND word251 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2082 Y0 word310 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2083 GND word465 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2084 Y6 word406 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2085 GND word751 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2086 GND word367 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2087 Y4 word206 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2088 GND word697 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2089 Y4 word694 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2090 GND word335 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2091 Y4 word142 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2092 Y0 word292 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2093 Y5 word454 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2094 Y1 word604 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2095 Y0 word622 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2096 Y2 word900 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2097 Y6 word924 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2098 GND word865 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2099 GND word169 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2100 GND word229 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2101 GND word559 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2102 Y2 word166 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2103 GND word1005 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2104 Y2 word734 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2105 GND word157 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2106 Y5 word278 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2107 Y7 word376 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2108 Y2 word654 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2109 Y6 word970 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2110 GND word495 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2111 GND word783 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2112 Y1 word484 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2113 Y2 word1000 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2114 Y6 word748 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2115 GND word271 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2116 GND word839 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X2117 GND word151 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2118 Y1 word262 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2119 GND word429 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2120 GND word203 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2121 Y7 word422 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2122 Y3 word888 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2123 Y7 word358 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2124 Y1 word528 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2125 Y2 word534 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2126 Y7 word688 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2127 GND word375 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2128 GND word253 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2129 Y2 word312 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2130 Y5 word480 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2131 GND word417 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X2132 GND word575 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2133 GND word687 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2134 Y2 word192 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2135 Y3 word504 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2136 Y1 word740 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2137 Y2 word680 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2138 Y6 word164 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2139 GND word915 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X2140 Y0 word974 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2141 GND word947 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2142 GND word851 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X2143 Y0 word216 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2144 GND word371 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2145 Y5 word940 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2146 Y6 word210 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2147 Y3 word328 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2148 Y7 word716 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2149 Y3 word384 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2150 Y4 word952 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2151 GND word893 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2152 Y6 word146 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2153 GND word171 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2154 GND word321 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2155 Y6 word476 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2156 GND word1015 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X2157 Y3 word162 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2158 Y1 word988 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2159 GND word659 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2160 GND word591 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2161 Y3 word650 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2162 Y4 word378 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2163 GND word489 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2164 Y5 word922 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2165 GND word727 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2166 GND word155 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2167 GND word251 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2168 Y6 word310 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2169 Y4 word434 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2170 Y3 word208 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2171 GND word425 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2172 Y0 word584 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2173 GND word153 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2174 Y4 word212 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2175 Y0 word362 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2176 GND word483 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2177 GND word201 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2178 Y7 word862 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2179 GND word539 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2180 GND word935 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2181 Y1 word868 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X2182 GND word809 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2183 Y6 word292 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2184 GND word317 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2185 Y0 word408 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2186 GND word467 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2187 Y6 word622 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2188 Y7 word908 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2189 Y2 word804 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2190 Y6 word710 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2191 Y1 word224 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2192 Y0 word242 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2193 Y7 word742 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2194 GND word221 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2195 Y6 word874 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2196 GND word815 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2197 Y0 word508 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2198 GND word179 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2199 GND word845 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2200 Y2 word786 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2201 Y7 word428 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2202 GND word955 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X2203 Y7 word326 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2204 GND word979 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2205 Y5 word386 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2206 GND word595 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2207 GND word733 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2208 GND word891 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2209 Y6 word856 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2210 Y3 word730 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2211 GND word161 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2212 Y5 word220 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2213 GND word379 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2214 Y1 word370 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2215 GND word491 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2216 Y5 word550 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2217 Y1 word700 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2218 GND word157 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2219 Y3 word996 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2220 Y1 word148 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2221 GND word367 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2222 GND word427 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2223 GND word645 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2224 GND word961 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2225 GND word697 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2226 Y7 word206 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2227 Y2 word484 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X2228 Y1 word636 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2229 Y7 word694 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2230 Y7 word142 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2231 GND word203 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2232 GND word413 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2233 Y0 word714 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2234 Y2 word528 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2235 GND word525 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2236 Y0 word760 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2237 GND word303 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2238 Y6 word216 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2239 GND word573 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2240 Y2 word630 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2241 GND word229 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2242 GND word897 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2243 Y0 word166 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2244 GND word559 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2245 GND word797 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2246 Y1 word894 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2247 Y5 word890 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2248 Y4 word794 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2249 Y3 word278 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2250 Y0 word654 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2251 GND word155 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2252 Y3 word334 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2253 Y4 word902 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2254 GND word271 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2255 GND word429 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2256 Y0 word906 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2257 Y6 word584 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2258 GND word929 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2259 GND word899 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2260 GND word541 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2261 Y5 word872 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2262 Y6 word362 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2263 Y0 word478 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2264 GND word707 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2265 GND word201 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2266 Y4 word384 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2267 GND word633 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2268 GND word375 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2269 Y0 word534 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2270 Y4 word162 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2271 GND word253 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2272 Y0 word312 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2273 Y6 word408 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2274 GND word467 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2275 GND word753 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2276 GND word885 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2277 Y3 word480 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2278 Y0 word578 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2279 Y4 word208 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2280 Y6 word242 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2281 GND word417 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2282 Y0 word634 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2283 GND word719 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2284 Y4 word696 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2285 GND word353 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2286 GND word687 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2287 Y1 word174 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2288 GND word853 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2289 Y0 word192 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2290 Y4 word530 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2291 Y6 word926 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2292 GND word859 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2293 GND word171 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2294 Y6 word824 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2295 Y0 word680 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2296 GND word231 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2297 Y1 word440 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2298 GND word765 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2299 GND word129 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2300 Y0 word458 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2301 GND word613 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2302 GND word659 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2303 Y7 word958 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2304 Y2 word736 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2305 Y2 word224 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2306 Y7 word378 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2307 GND word905 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2308 GND word215 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2309 GND word395 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2310 Y7 word434 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2311 GND word647 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2312 GND word153 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2313 Y7 word212 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2314 GND word999 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2315 Y5 word170 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2316 Y2 word718 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2317 Y1 word320 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2318 Y3 word946 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2319 GND word887 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2320 GND word377 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2321 GND word911 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2322 GND word527 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2323 GND word275 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2324 GND word823 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2325 Y2 word148 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2326 Y5 word482 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2327 Y1 word632 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2328 GND word691 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2329 Y1 word568 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2330 GND word923 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2331 Y1 word964 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2332 Y4 word864 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2333 Y6 word166 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2334 Y0 word976 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2335 GND word739 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2336 GND word179 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2337 GND word1005 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X2338 Y4 word454 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2339 Y0 word604 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2340 Y3 word386 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2341 Y6 word478 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2342 GND word229 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2343 GND word379 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2344 Y3 word652 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2345 GND word161 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2346 Y3 word220 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2347 GND word879 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2348 GND word157 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2349 GND word491 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2350 GND word881 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2351 Y5 word822 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X2352 Y0 word792 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X2353 GND word253 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2354 Y6 word312 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2355 Y4 word436 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2356 Y4 word334 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2357 GND word427 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2358 GND word325 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2359 Y0 word484 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2360 Y6 word578 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2361 GND word203 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2362 Y0 word262 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2363 GND word541 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2364 Y4 word600 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2365 Y6 word634 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2366 Y7 word920 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2367 Y7 word762 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2368 GND word353 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2369 Y5 word140 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2370 Y0 word528 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2371 GND word761 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2372 Y6 word192 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2373 Y3 word704 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2374 GND word303 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2375 Y5 word968 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2376 Y6 word458 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2377 Y4 word480 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2378 GND word573 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2379 Y6 word876 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2380 Y0 word630 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2381 Y3 word750 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2382 GND word181 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2383 Y5 word240 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2384 Y1 word390 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2385 GND word847 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2386 Y2 word788 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2387 GND word957 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X2388 Y2 word174 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2389 Y7 word328 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2390 GND word981 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2391 GND word165 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2392 GND word345 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2393 Y7 word384 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2394 GND word917 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2395 GND word893 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2396 Y6 word858 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2397 Y3 word732 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2398 Y7 word162 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2399 Y2 word440 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2400 Y6 word756 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2401 Y5 word222 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2402 GND word279 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2403 Y1 word372 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2404 Y7 word650 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2405 Y1 word270 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2406 Y5 word552 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2407 Y3 word998 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2408 GND word727 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2409 GND word211 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2410 GND word549 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2411 GND word647 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2412 GND word963 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2413 GND word215 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2414 Y3 word896 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2415 GND word837 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X2416 Y7 word208 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2417 GND word425 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2418 Y1 word536 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2419 Y7 word696 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2420 Y2 word320 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2421 GND word809 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2422 Y0 word716 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2423 GND word527 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2424 GND word821 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2425 Y1 word914 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2426 Y5 word698 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2427 Y1 word850 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2428 Y2 word632 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2429 Y6 word604 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2430 GND word623 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2431 GND word231 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2432 Y2 word568 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2433 GND word129 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2434 Y0 word862 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2435 GND word955 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2436 Y0 word224 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2437 GND word379 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2438 Y4 word404 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2439 GND word497 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2440 Y0 word554 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2441 Y3 word336 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2442 GND word395 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2443 Y7 word724 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2444 GND word157 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2445 GND word901 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2446 GND word179 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2447 GND word329 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2448 Y3 word602 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2449 Y3 word170 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2450 Y1 word838 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2451 GND word989 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2452 GND word831 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X2453 Y0 word742 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2454 GND word203 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2455 Y4 word386 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2456 GND word161 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2457 Y4 word220 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2458 Y4 word942 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2459 GND word1001 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2460 Y0 word370 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2461 Y0 word700 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2462 Y3 word482 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2463 Y7 word870 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2464 Y0 word148 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2465 GND word303 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2466 Y0 word636 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2467 GND word475 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2468 GND word721 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2469 Y6 word630 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2470 GND word235 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2471 Y4 word532 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2472 Y6 word928 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2473 Y3 word802 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2474 Y0 word682 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2475 GND word523 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2476 Y6 word826 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2477 GND word767 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X2478 GND word131 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2479 Y5 word190 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2480 GND word229 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2481 Y1 word340 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2482 GND word797 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X2483 GND word619 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2484 Y3 word966 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2485 GND word907 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2486 GND word217 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2487 GND word397 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2488 Y7 word436 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2489 GND word547 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2490 Y7 word334 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2491 GND word573 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2492 Y2 word902 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2493 Y5 word394 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2494 GND word867 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2495 GND word899 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2496 Y5 word172 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2497 Y1 word322 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2498 GND word1007 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2499 GND word597 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2500 Y6 word972 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2501 GND word913 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2502 GND word165 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2503 Y1 word588 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2504 Y1 word156 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2505 GND word277 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2506 GND word375 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2507 Y1 word486 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2508 Y5 word494 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2509 Y1 word644 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2510 GND word213 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2511 Y2 word372 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2512 GND word211 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2513 GND word641 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2514 GND word759 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2515 Y2 word702 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2516 Y2 word638 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2517 Y3 word140 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2518 GND word477 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2519 Y2 word536 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2520 Y5 word318 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2521 Y1 word468 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2522 GND word929 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2523 GND word687 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2524 Y4 word764 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2525 GND word311 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2526 Y0 word978 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2527 GND word859 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X2528 GND word971 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2529 Y6 word224 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2530 Y3 word240 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2531 GND word181 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2532 Y2 word518 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2533 Y0 word812 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2534 Y0 word174 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2535 GND word805 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2536 GND word623 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2537 GND word231 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2538 GND word129 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2539 Y3 word222 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2540 Y0 word440 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2541 GND word595 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2542 Y4 word910 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2543 GND word279 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2544 Y7 word940 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2545 GND word497 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2546 Y1 word946 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X2547 GND word883 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2548 GND word215 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2549 GND word939 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X2550 Y5 word880 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2551 Y4 word336 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2552 Y6 word370 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2553 GND word715 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2554 GND word327 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2555 Y6 word148 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2556 Y4 word170 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2557 GND word577 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2558 Y4 word602 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2559 Y6 word636 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2560 Y7 word922 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2561 GND word951 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2562 Y4 word892 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2563 Y0 word320 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2564 GND word475 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2565 GND word649 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2566 GND word377 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2567 GND word763 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2568 Y3 word368 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2569 Y0 word586 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2570 Y3 word698 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2571 GND word185 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2572 GND word361 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2573 Y7 word404 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2574 Y4 word482 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2575 Y0 word632 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2576 Y6 word878 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2577 GND word861 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2578 Y3 word752 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2579 GND word473 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2580 Y6 word934 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2581 GND word969 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2582 GND word179 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2583 GND word239 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2584 Y0 word568 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2585 Y6 word712 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2586 GND word235 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2587 Y1 word226 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2588 GND word445 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2589 Y2 word744 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2590 GND word167 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2591 GND word347 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2592 Y7 word386 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2593 Y5 word564 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2594 Y3 word852 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2595 GND word283 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2596 Y5 word344 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2597 Y2 word1010 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X2598 GND word817 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2599 Y6 word758 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2600 GND word161 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2601 Y7 word220 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2602 Y2 word340 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2603 Y7 word652 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2604 Y1 word272 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2605 GND word217 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2606 Y5 word610 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2607 Y3 word898 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2608 GND word427 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2609 Y5 word388 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2610 GND word325 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2611 Y2 word992 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X2612 GND word163 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2613 Y2 word156 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2614 Y1 word704 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2615 GND word699 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2616 Y1 word418 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2617 GND word363 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2618 GND word693 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2619 Y4 word140 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2620 Y6 word174 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2621 Y0 word984 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2622 GND word131 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2623 Y3 word190 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2624 Y2 word468 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X2625 Y4 word916 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2626 Y1 word1016 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2627 Y0 word762 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2628 GND word285 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2629 GND word619 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2630 GND word755 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2631 Y3 word394 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2632 Y1 word732 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2633 GND word181 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2634 GND word215 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2635 Y4 word240 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2636 Y0 word390 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2637 Y4 word962 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2638 Y3 word172 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2639 Y7 word890 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2640 GND word991 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2641 Y1 word896 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2642 GND word837 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X2643 Y4 word796 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2644 GND word165 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2645 GND word345 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2646 GND word889 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2647 Y5 word830 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2648 Y6 word320 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2649 GND word277 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2650 GND word1003 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2651 Y4 word222 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2652 Y0 word372 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2653 GND word431 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2654 GND word213 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2655 Y6 word586 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2656 GND word931 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2657 Y7 word872 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2658 Y4 word842 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2659 GND word709 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2660 Y0 word702 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2661 GND word211 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2662 Y0 word270 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2663 GND word543 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2664 Y0 word638 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2665 GND word309 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2666 GND word361 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2667 Y3 word318 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2668 GND word477 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2669 Y0 word536 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2670 Y6 word632 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2671 Y7 word706 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2672 GND word593 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2673 GND word135 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2674 GND word311 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2675 GND word919 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2676 Y6 word828 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2677 GND word231 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2678 Y6 word884 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2679 GND word129 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2680 GND word133 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2681 Y4 word368 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2682 Y0 word518 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2683 GND word189 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2684 GND word855 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2685 Y4 word698 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2686 GND word185 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2687 Y1 word176 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2688 GND word395 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2689 Y7 word336 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2690 GND word455 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2691 Y1 word664 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2692 GND word233 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2693 GND word925 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2694 GND word901 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2695 Y7 word170 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2696 Y5 word230 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2697 Y1 word380 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2698 GND word167 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2699 Y2 word226 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2700 Y5 word560 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2701 Y3 word1006 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2702 Y1 word158 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2703 GND word377 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2704 Y5 word338 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2705 Y1 word488 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2706 GND word433 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X2707 Y2 word942 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X2708 GND word1001 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2709 GND word331 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X2710 Y1 word544 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2711 GND word643 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2712 Y2 word272 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2713 Y0 word724 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2714 Y4 word766 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2715 Y3 word464 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2716 Y1 word802 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X2717 GND word239 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2718 GND word907 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2719 Y4 word866 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2720 GND word807 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2721 GND word235 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2722 Y6 word390 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2723 Y5 word900 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2724 GND word735 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2725 GND word505 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2726 Y3 word344 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2727 GND word131 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2728 GND word165 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2729 Y4 word190 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2730 GND word281 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2731 Y0 word340 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2732 GND word597 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2733 Y4 word912 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2734 Y7 word840 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2735 GND word1007 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X2736 Y4 word848 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2737 GND word669 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2738 GND word217 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2739 Y6 word372 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2740 GND word941 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2741 GND word717 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2742 GND word211 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2743 Y1 word782 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2744 GND word723 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2745 Y5 word154 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2746 Y6 word638 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2747 GND word953 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2748 Y4 word172 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2749 Y0 word322 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2750 GND word381 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2751 GND word163 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2752 GND word477 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2753 GND word881 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2754 Y4 word660 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2755 GND word651 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2756 Y7 word140 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2757 Y4 word438 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2758 Y0 word588 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2759 Y0 word156 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2760 GND word311 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2761 Y0 word486 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2762 Y0 word644 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2763 GND word729 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2764 GND word213 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2765 GND word363 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2766 GND word543 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2767 GND word261 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2768 GND word863 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2769 GND word599 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2770 Y6 word936 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2771 GND word971 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X2772 GND word761 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2773 GND word181 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2774 Y7 word240 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2775 Y4 word318 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2776 Y1 word450 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2777 Y0 word468 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2778 GND word139 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2779 GND word623 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2780 GND word135 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2781 Y1 word228 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2782 GND word447 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2783 GND word711 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2784 GND word345 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2785 Y5 word566 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2786 GND word225 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2787 Y1 word284 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2788 Y2 word1012 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2789 GND word555 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2790 GND word851 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2791 GND word183 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2792 Y7 word222 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2793 GND word875 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2794 GND word749 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2795 Y5 word612 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2796 Y5 word180 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2797 Y1 word330 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2798 GND word787 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2799 Y2 word176 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2800 Y3 word956 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2801 GND word327 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2802 GND word605 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2803 Y6 word980 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2804 Y2 word664 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2805 GND word387 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2806 Y1 word596 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2807 GND word655 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2808 GND word383 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2809 Y2 word892 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2810 Y2 word380 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2811 Y1 word430 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2812 Y5 word492 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2813 GND word551 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2814 GND word649 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2815 Y2 word158 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2816 GND word309 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2817 Y7 word368 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2818 Y2 word488 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2819 Y2 word646 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2820 Y2 word544 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2821 Y7 word698 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2822 GND word263 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2823 Y5 word804 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X2824 Y1 word752 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2825 GND word235 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2826 GND word745 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2827 GND word133 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2828 GND word189 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2829 GND word757 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2830 GND word185 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2831 GND word909 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2832 Y4 word464 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X2833 GND word793 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2834 GND word845 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2835 GND word217 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2836 GND word849 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X2837 GND word233 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2838 GND word239 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2839 Y3 word230 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2840 Y3 word560 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2841 Y1 word898 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2842 GND word861 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X2843 GND word167 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2844 Y0 word226 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2845 GND word347 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2846 GND word381 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2847 Y4 word564 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2848 GND word891 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2849 Y3 word496 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2850 Y7 word726 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2851 GND word283 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2852 GND word433 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2853 Y6 word588 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2854 GND word903 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2855 Y6 word156 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2856 Y0 word272 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2857 GND word331 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2858 GND word933 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2859 GND word669 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2860 Y3 word542 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2861 GND word601 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2862 Y6 word904 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2863 GND word363 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2864 Y4 word388 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2865 Y0 word538 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2866 GND word873 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2867 Y7 word708 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2868 GND word209 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2869 Y2 word816 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2870 Y0 word594 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2871 Y3 word714 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2872 GND word145 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2873 GND word163 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2874 Y1 word354 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2875 GND word313 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2876 Y6 word468 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2877 GND word921 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2878 Y6 word886 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2879 GND word819 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2880 GND word131 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2881 Y7 word190 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2882 Y5 word250 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2883 Y4 word268 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2884 Y1 word400 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2885 Y0 word418 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2886 Y6 word720 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2887 Y1 word178 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2888 GND word397 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2889 Y1 word234 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2890 GND word457 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2891 GND word175 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2892 Y7 word394 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2893 GND word927 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2894 GND word509 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2895 GND word801 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2896 Y7 word172 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2897 Y5 word232 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2898 GND word825 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2899 Y1 word500 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2900 Y5 word562 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2901 GND word621 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2902 Y7 word660 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2903 Y5 word130 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2904 Y2 word228 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2905 Y1 word280 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2906 Y2 word796 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2907 GND word225 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2908 Y2 word284 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X2909 Y7 word438 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2910 Y3 word906 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2911 Y2 word614 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2912 GND word337 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2913 Y5 word396 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2914 Y3 word154 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2915 GND word213 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2916 Y2 word842 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2917 GND word785 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2918 GND word389 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2919 GND word655 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2920 GND word587 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2921 GND word919 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2922 Y5 word754 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2923 GND word701 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2924 GND word185 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2925 Y1 word692 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2926 GND word359 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2927 GND word637 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2928 GND word931 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2929 GND word139 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2930 GND word865 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2931 GND word135 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2932 GND word743 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2933 Y6 word226 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2934 Y0 word706 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2935 GND word133 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2936 GND word167 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2937 GND word799 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X2938 GND word183 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2939 GND word189 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2940 Y3 word180 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2941 GND word943 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2942 GND word671 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2943 Y0 word176 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2944 GND word811 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2945 GND word455 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X2946 GND word387 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2947 Y0 word664 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2948 GND word233 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2949 Y0 word1018 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X2950 GND word383 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2951 Y4 word230 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2952 Y0 word380 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2953 GND word439 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2954 GND word883 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2955 Y6 word594 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2956 GND word653 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2957 GND word939 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2958 Y7 word880 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2959 Y0 word158 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2960 Y5 word882 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2961 GND word313 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2962 Y0 word488 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X2963 Y4 word496 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X2964 Y0 word646 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X2965 GND word823 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2966 Y2 word766 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2967 GND word731 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2968 Y0 word544 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X2969 GND word245 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2970 Y1 word304 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2971 GND word263 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X2972 GND word601 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2973 Y4 word542 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2974 Y3 word592 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2975 GND word895 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2976 GND word871 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X2977 GND word763 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2978 GND word923 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2979 Y5 word200 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2980 GND word239 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2981 Y2 word866 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2982 Y1 word350 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2983 GND word807 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X2984 GND word295 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X2985 Y3 word976 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2986 Y1 word128 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2987 Y1 word286 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X2988 GND word347 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X2989 Y1 word184 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2990 Y1 word616 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2991 Y7 word344 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2992 Y2 word912 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X2993 GND word877 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2994 Y3 word810 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X2995 GND word751 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2996 Y5 word182 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X2997 GND word241 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X2998 Y2 word400 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X2999 GND word669 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3000 Y2 word178 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3001 GND word175 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3002 Y2 word234 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3003 Y7 word388 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3004 Y5 word448 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3005 Y7 word444 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3006 Y5 word346 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3007 Y6 word918 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3008 GND word953 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X3009 GND word163 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3010 GND word441 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3011 Y2 word500 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3012 GND word223 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3013 Y5 word282 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3014 GND word339 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X3015 Y1 word432 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3016 GND word651 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3017 Y2 word280 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3018 GND word553 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3019 GND word703 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3020 GND word209 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3021 Y4 word154 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3022 GND word145 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3023 GND word135 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3024 Y3 word250 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3025 Y0 word822 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X3026 GND word457 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3027 GND word847 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3028 Y6 word176 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3029 Y4 word300 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3030 Y0 word450 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3031 GND word509 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3032 GND word139 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3033 Y3 word232 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3034 GND word605 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3035 Y7 word950 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3036 Y3 word130 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3037 Y0 word228 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3038 GND word621 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3039 GND word893 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3040 GND word863 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3041 GND word383 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3042 Y4 word566 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3043 GND word1015 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X3044 Y7 word728 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3045 GND word225 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3046 Y0 word284 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3047 Y6 word380 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3048 GND word405 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3049 Y3 word498 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3050 Y0 word614 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3051 GND word949 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3052 GND word725 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3053 Y6 word158 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3054 GND word183 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3055 Y0 word968 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3056 GND word333 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3057 GND word961 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X3058 GND word671 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3059 Y4 word180 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3060 Y0 word330 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3061 GND word389 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3062 GND word603 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3063 GND word833 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3064 GND word993 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3065 GND word889 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3066 GND word387 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3067 Y0 word596 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3068 Y3 word716 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3069 Y6 word740 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3070 GND word147 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3071 GND word195 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3072 Y1 word254 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3073 Y7 word414 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3074 Y0 word430 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3075 GND word133 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3076 Y7 word930 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3077 GND word821 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3078 Y5 word252 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3079 GND word189 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3080 GND word757 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X3081 Y6 word722 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3082 GND word245 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3083 Y2 word304 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3084 Y1 word236 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3085 Y5 word416 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3086 Y1 word134 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3087 Y5 word574 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3088 GND word233 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3089 GND word827 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3090 Y5 word352 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3091 GND word409 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3092 Y1 word502 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3093 Y5 word132 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3094 GND word191 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3095 Y7 word230 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3096 Y2 word128 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3097 GND word679 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3098 Y7 word338 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3099 Y2 word616 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3100 GND word967 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X3101 Y3 word908 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3102 Y2 word184 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3103 Y1 word218 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3104 Y5 word398 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3105 Y1 word548 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3106 GND word607 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3107 GND word903 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3108 Y6 word868 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3109 GND word173 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3110 Y1 word382 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3111 Y3 word1008 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3112 Y2 word598 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3113 GND word973 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3114 Y1 word648 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3115 GND word985 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X3116 GND word885 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3117 Y2 word432 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3118 Y0 word726 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3119 Y7 word642 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3120 GND word703 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3121 Y1 word760 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3122 GND word209 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3123 Y3 word302 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3124 Y3 word200 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3125 GND word145 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3126 Y0 word354 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3127 Y4 word926 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3128 Y0 word772 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3129 GND word295 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3130 Y6 word450 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3131 Y7 word854 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3132 GND word765 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3133 Y3 word466 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3134 Y0 word708 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3135 Y6 word228 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3136 Y5 word738 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3137 GND word225 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3138 Y4 word250 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3139 Y0 word400 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3140 GND word459 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3141 Y6 word614 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3142 Y3 word182 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3143 GND word241 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3144 GND word959 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3145 Y7 word900 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3146 Y0 word178 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3147 Y5 word902 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3148 GND word843 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3149 Y1 word906 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3150 Y4 word806 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3151 Y0 word666 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3152 GND word175 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3153 Y0 word234 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3154 GND word389 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3155 Y3 word448 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3156 GND word507 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3157 GND word899 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3158 Y7 word154 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3159 Y7 word734 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3160 Y4 word232 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3161 GND word441 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3162 Y0 word500 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3163 Y4 word562 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3164 Y6 word596 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3165 GND word911 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3166 Y4 word130 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3167 GND word223 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3168 Y0 word280 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3169 GND word339 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3170 GND word553 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3171 GND word941 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3172 GND word839 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3173 Y4 word498 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3174 Y0 word546 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3175 Y1 word204 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3176 GND word603 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3177 GND word637 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3178 Y4 word662 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3179 GND word897 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3180 GND word359 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3181 Y5 word202 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3182 GND word437 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3183 Y6 word894 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3184 GND word139 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3185 Y3 word978 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3186 GND word865 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3187 GND word195 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3188 Y2 word254 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3189 Y1 word288 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3190 Y1 word186 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3191 GND word405 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3192 Y6 word938 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3193 Y0 word692 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3194 GND word183 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3195 GND word243 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3196 Y1 word452 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3197 GND word671 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3198 Y7 word180 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3199 GND word713 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3200 GND word629 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3201 Y2 word236 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3202 Y2 word134 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3203 Y1 word168 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3204 GND word227 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3205 Y5 word348 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3206 GND word387 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3207 Y7 word446 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3208 GND word565 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3209 GND word853 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3210 GND word1011 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3211 Y6 word818 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3212 GND word653 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3213 Y1 word332 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3214 GND word611 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3215 Y2 word218 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3216 GND word607 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3217 GND word147 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3218 GND word323 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X3219 Y6 word354 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3220 GND word295 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3221 Y3 word252 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3222 Y2 word648 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3223 GND word883 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X3224 Y0 word304 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3225 Y1 word976 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3226 Y0 word880 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3227 Y4 word876 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3228 GND word245 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3229 Y6 word400 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3230 GND word459 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3231 GND word969 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3232 Y3 word416 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3233 Y3 word574 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3234 GND word745 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3235 Y6 word178 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3236 Y4 word302 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3237 Y1 word810 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3238 GND word751 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3239 GND word747 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3240 Y4 word200 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3241 Y6 word234 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3242 GND word293 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3243 Y3 word352 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3244 Y5 word744 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3245 GND word175 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3246 Y0 word350 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3247 GND word409 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3248 Y3 word132 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3249 GND word191 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3250 GND word1017 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3251 GND word909 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3252 Y0 word128 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3253 Y0 word286 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3254 Y0 word184 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3255 GND word407 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3256 Y4 word466 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3257 Y0 word616 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3258 GND word845 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3259 Y4 word756 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3260 Y4 word182 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3261 GND word241 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3262 GND word963 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3263 GND word173 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3264 GND word391 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3265 GND word891 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3266 Y4 word448 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3267 Y6 word964 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3268 Y5 word992 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3269 GND word209 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3270 Y0 word598 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3271 Y4 word346 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3272 GND word145 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3273 GND word739 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3274 GND word223 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3275 Y4 word282 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3276 Y0 word432 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3277 GND word373 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3278 GND word587 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3279 Y7 word932 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3280 Y2 word710 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3281 GND word873 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3282 Y7 word250 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3283 GND word369 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3284 GND word519 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3285 Y2 word874 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3286 GND word815 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3287 Y2 word204 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3288 Y1 word238 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3289 Y5 word576 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3290 GND word635 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3291 Y3 word984 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3292 Y1 word136 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3293 Y5 word144 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3294 Y1 word294 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3295 Y1 word624 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3296 Y3 word920 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3297 Y6 word888 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3298 Y3 word762 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3299 Y7 word232 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3300 GND word979 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X3301 GND word193 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3302 Y1 word402 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3303 Y7 word130 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3304 GND word249 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3305 Y2 word288 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3306 Y2 word856 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3307 GND word681 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3308 Y2 word186 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3309 GND word177 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3310 GND word337 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3311 Y7 word396 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3312 Y5 word456 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3313 GND word803 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3314 GND word393 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3315 Y2 word452 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3316 GND word961 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X3317 GND word449 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3318 Y7 word662 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3319 Y2 word168 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3320 GND word227 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3321 GND word561 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3322 Y5 word620 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3323 GND word437 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3324 GND word557 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3325 Y1 word716 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3326 GND word1009 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3327 GND word493 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3328 Y0 word728 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3329 Y2 word332 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3330 GND word721 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X3331 GND word245 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3332 Y6 word304 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3333 Y3 word202 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3334 Y4 word928 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3335 GND word833 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X3336 GND word147 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3337 GND word195 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3338 Y0 word254 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3339 GND word889 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3340 Y0 word830 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X3341 GND word767 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3342 GND word409 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3343 Y7 word754 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3344 Y3 word524 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3345 Y6 word128 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3346 Y4 word252 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3347 Y6 word184 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3348 GND word243 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3349 Y6 word616 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3350 GND word967 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3351 Y1 word908 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3352 Y4 word808 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3353 Y0 word236 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3354 Y4 word416 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3355 Y0 word930 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3356 GND word901 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3357 Y0 word134 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3358 GND word391 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3359 Y4 word574 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3360 Y7 word736 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3361 Y3 word506 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3362 Y4 word352 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3363 GND word443 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3364 Y0 word502 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3365 Y4 word132 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3366 GND word191 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3367 Y6 word598 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3368 GND word943 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3369 Y4 word972 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3370 GND word913 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3371 GND word341 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3372 GND word499 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3373 Y1 word1008 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3374 Y6 word914 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3375 GND word841 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3376 Y3 word670 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3377 Y0 word218 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3378 GND word373 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3379 Y5 word942 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3380 Y0 word548 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3381 Y7 word718 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3382 GND word173 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3383 Y5 word214 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3384 GND word323 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3385 Y1 word364 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3386 Y0 word382 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3387 GND word485 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3388 Y3 word990 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3389 Y7 word882 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3390 GND word719 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3391 GND word661 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3392 Y7 word200 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3393 Y0 word648 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3394 GND word319 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3395 Y2 word926 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3396 GND word733 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3397 GND word487 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3398 Y2 word824 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3399 GND word247 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3400 GND word765 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3401 Y6 word730 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3402 Y1 word188 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3403 GND word407 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3404 GND word423 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3405 Y1 word244 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3406 GND word923 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3407 Y7 word182 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3408 GND word241 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3409 GND word519 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3410 Y1 word510 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3411 Y5 word690 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3412 GND word199 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3413 Y2 word238 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3414 GND word631 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3415 Y2 word806 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3416 Y2 word136 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3417 Y7 word346 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3418 GND word567 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3419 Y2 word624 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3420 GND word1013 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3421 Y1 word556 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3422 GND word615 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3423 GND word223 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3424 GND word343 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3425 GND word911 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3426 Y0 word854 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X3427 GND word795 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3428 GND word177 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3429 Y1 word656 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3430 GND word959 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3431 GND word929 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3432 Y0 word734 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3433 GND word195 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3434 Y6 word254 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3435 Y5 word764 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3436 GND word707 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3437 Y4 word878 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3438 GND word941 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X3439 Y0 word1000 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X3440 Y0 word204 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3441 GND word839 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X3442 Y3 word144 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3443 Y3 word576 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3444 GND word635 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3445 Y3 word474 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3446 Y1 word812 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3447 Y4 word202 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3448 Y6 word236 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3449 GND word983 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3450 GND word805 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3451 Y5 word746 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3452 Y6 word134 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3453 GND word193 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3454 GND word681 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3455 GND word249 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3456 Y0 word288 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3457 GND word817 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X3458 Y4 word758 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3459 Y0 word186 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3460 Y5 word910 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3461 GND word847 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3462 GND word853 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.2193 ps=1.88 w=0.51 l=0.17
X3463 Y0 word674 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3464 Y3 word456 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3465 Y5 word846 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3466 GND word759 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3467 Y6 word218 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3468 GND word243 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3469 GND word393 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3470 Y0 word452 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3471 GND word299 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3472 GND word607 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3473 Y7 word952 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3474 GND word893 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3475 GND word449 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3476 GND word629 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3477 Y3 word620 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3478 GND word949 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3479 Y1 word958 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X3480 Y0 word168 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3481 GND word227 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3482 Y4 word348 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3483 Y6 word382 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3484 GND word565 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3485 Y5 word892 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3486 GND word859 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3487 GND word727 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3488 GND word147 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3489 Y5 word164 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3490 GND word493 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3491 GND word273 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3492 Y1 word314 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3493 Y0 word332 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3494 Y3 word940 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3495 Y7 word832 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3496 Y4 word670 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3497 Y7 word252 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3498 GND word905 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3499 GND word371 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3500 Y5 word210 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3501 GND word715 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3502 Y1 word138 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3503 Y5 word146 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3504 GND word197 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3505 Y2 word364 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3506 Y7 word416 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3507 Y1 word194 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3508 Y7 word352 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3509 GND word887 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3510 Y3 word820 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3511 Y7 word132 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3512 GND word191 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3513 GND word469 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3514 GND word251 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3515 Y5 word310 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3516 Y1 word460 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3517 GND word917 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X3518 GND word679 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3519 Y2 word188 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3520 GND word247 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3521 Y7 word398 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3522 Y2 word244 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3523 GND word667 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3524 GND word963 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X3525 GND word173 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3526 Y0 word804 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3527 Y1 word442 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3528 GND word563 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3529 Y5 word622 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3530 GND word661 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3531 GND word615 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3532 GND word909 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X3533 Y3 word214 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3534 GND word845 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3535 Y6 word204 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3536 GND word319 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3537 Y2 word656 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3538 Y4 word828 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3539 VDD GND Y6 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X3540 Y4 word884 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3541 Y3 word526 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3542 GND word585 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3543 Y5 word916 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3544 Y1 word920 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X3545 Y6 word186 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3546 GND word755 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3547 GND word301 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3548 Y3 word360 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3549 GND word873 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3550 GND word199 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3551 Y0 word238 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3552 GND word297 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3553 GND word393 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3554 Y6 word452 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3555 Y4 word576 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3556 GND word635 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3557 Y5 word962 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3558 Y0 word136 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3559 Y4 word144 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3560 Y0 word294 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3561 Y7 word738 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3562 GND word449 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3563 Y0 word624 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3564 GND word465 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3565 GND word737 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3566 Y6 word168 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3567 GND word193 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3568 GND word227 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3569 GND word343 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3570 Y0 word402 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3571 GND word249 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3572 Y7 word902 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3573 GND word843 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3574 GND word399 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3575 Y3 word672 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3576 GND word159 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3577 GND word899 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3578 GND word177 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3579 GND word785 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3580 Y5 word216 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3581 Y6 word750 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3582 Y1 word264 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3583 GND word561 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3584 Y3 word890 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3585 Y7 word202 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3586 Y2 word826 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3587 GND word767 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3588 Y6 word732 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3589 GND word155 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3590 Y1 word246 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3591 Y3 word872 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3592 GND word243 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3593 Y6 word896 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3594 GND word571 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3595 GND word633 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3596 GND word201 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3597 Y1 word410 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3598 Y2 word138 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3599 GND word197 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3600 GND word355 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X3601 GND word977 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3602 GND word689 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3603 Y7 word348 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3604 GND word685 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3605 Y2 word194 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3606 Y1 word676 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3607 GND word937 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3608 GND word913 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3609 Y5 word242 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3610 GND word401 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3611 Y2 word460 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3612 Y0 word754 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3613 Y1 word392 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3614 Y7 word670 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3615 Y4 word954 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X3616 Y1 word724 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3617 Y3 word164 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3618 GND word501 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3619 Y1 word990 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X3620 Y5 word766 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3621 Y0 word736 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3622 GND word613 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3623 GND word829 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X3624 GND word729 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3625 GND word269 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3626 GND word943 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3627 Y3 word210 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3628 Y2 word606 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3629 GND word995 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3630 GND word841 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X3631 Y4 word214 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3632 Y0 word364 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3633 GND word999 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3634 Y3 word146 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3635 GND word485 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3636 Y7 word864 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3637 GND word297 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3638 GND word807 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3639 GND word777 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3640 Y0 word718 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3641 Y6 word238 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3642 Y1 word870 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X3643 Y6 word136 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3644 Y6 word294 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3645 GND word319 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3646 GND word469 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3647 GND word251 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3648 Y3 word310 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3649 Y6 word624 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3650 GND word247 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3651 Y0 word188 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3652 Y6 word402 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3653 GND word975 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3654 Y5 word912 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3655 GND word747 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3656 Y0 word244 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3657 GND word399 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3658 Y5 word848 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3659 Y7 word744 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3660 GND word177 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3661 GND word301 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3662 Y0 word510 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3663 GND word199 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3664 GND word631 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3665 Y4 word690 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3666 GND word349 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3667 Y3 word622 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3668 GND word567 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3669 Y4 word406 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3670 GND word465 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3671 GND word735 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3672 Y0 word556 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3673 Y5 word166 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3674 Y1 word316 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3675 Y4 word672 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3676 Y6 word966 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3677 GND word159 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3678 GND word907 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3679 Y3 word840 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3680 Y1 word150 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3681 GND word369 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3682 GND word429 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3683 Y0 word656 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3684 GND word717 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3685 GND word741 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3686 Y2 word264 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3687 Y7 word144 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3688 GND word255 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3689 Y2 word712 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3690 Y1 word196 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3691 GND word415 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3692 GND word193 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3693 GND word253 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3694 Y5 word312 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3695 GND word249 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3696 Y1 word462 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3697 GND word681 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3698 Y2 word758 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3699 GND word723 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3700 Y2 word246 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3701 GND word237 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3702 Y1 word296 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3703 GND word417 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3704 GND word575 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3705 Y5 word634 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3706 GND word761 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3707 Y5 word192 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3708 GND word351 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3709 GND word683 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3710 Y1 word342 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3711 Y5 word680 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3712 GND word287 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3713 Y5 word458 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3714 Y1 word608 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3715 Y4 word904 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3716 Y3 word216 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3717 Y2 word392 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3718 GND word847 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X3719 Y0 word788 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3720 Y6 word364 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3721 GND word709 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3722 GND word893 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3723 GND word715 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3724 Y4 word886 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3725 Y4 word164 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3726 Y0 word314 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3727 GND word469 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3728 GND word155 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3729 Y1 word922 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X3730 GND word247 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3731 GND word757 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3732 Y6 word188 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3733 Y1 word820 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3734 Y4 word210 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3735 Y6 word244 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3736 GND word269 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3737 GND word419 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3738 GND word201 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3739 GND word633 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3740 GND word993 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3741 Y0 word138 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3742 Y4 word146 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3743 GND word197 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3744 GND word927 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3745 Y4 word986 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3746 GND word773 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3747 GND word355 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3748 GND word535 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3749 Y0 word194 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3750 Y3 word408 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3751 GND word467 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3752 Y0 word626 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3753 GND word855 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3754 GND word861 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X3755 Y5 word798 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3756 GND word251 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3757 GND word401 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3758 Y0 word460 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3759 Y3 word242 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3760 GND word615 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3761 Y7 word960 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3762 GND word901 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3763 GND word903 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3764 Y2 word1004 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3765 Y6 word752 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3766 Y7 word214 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3767 Y1 word266 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3768 Y0 word442 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3769 GND word501 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3770 GND word563 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3771 Y7 word942 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3772 GND word779 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3773 GND word379 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3774 Y0 word606 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3775 Y2 word316 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3776 GND word157 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3777 Y1 word366 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3778 GND word205 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3779 GND word933 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X3780 GND word663 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3781 Y5 word484 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3782 Y6 word898 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3783 GND word831 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3784 Y2 word150 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3785 GND word421 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3786 GND word989 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3787 GND word141 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3788 GND word203 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3789 Y7 word360 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3790 Y1 word412 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3791 Y7 word690 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3792 GND word199 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3793 Y2 word196 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3794 GND word255 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3795 GND word187 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3796 Y7 word406 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3797 GND word675 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3798 Y7 word672 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3799 Y5 word630 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3800 GND word237 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3801 Y2 word296 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3802 GND word785 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3803 GND word1019 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3804 Y3 word166 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3805 GND word797 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3806 Y3 word654 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3807 Y1 word890 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3808 Y0 word738 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3809 GND word159 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3810 Y0 word794 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3811 Y4 word790 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3812 GND word731 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3813 Y6 word314 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3814 GND word271 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3815 Y2 word608 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3816 Y4 word216 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3817 GND word997 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3818 GND word895 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3819 Y0 word264 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3820 GND word899 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3821 GND word931 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X3822 Y1 word872 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X3823 Y7 word764 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3824 Y6 word138 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3825 GND word197 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3826 Y5 word924 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3827 GND word355 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3828 GND word471 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3829 Y6 word626 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3830 Y6 word194 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3831 GND word253 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3832 Y3 word312 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3833 GND word155 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3834 GND word877 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3835 Y0 word246 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3836 GND word305 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3837 GND word401 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3838 Y6 word460 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3839 Y5 word970 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3840 GND word417 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3841 GND word575 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3842 Y3 word634 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3843 Y7 word746 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3844 Y4 word362 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3845 Y5 word748 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3846 GND word633 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3847 Y4 word982 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X3848 GND word201 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3849 GND word351 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3850 Y0 word410 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3851 GND word683 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3852 Y3 word192 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3853 Y7 word910 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3854 GND word689 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3855 GND word287 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3856 GND word467 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3857 Y7 word846 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3858 Y0 word676 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3859 Y3 word458 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3860 GND word919 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3861 Y7 word164 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3862 Y5 word224 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3863 Y4 word242 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3864 Y0 word392 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3865 GND word451 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3866 Y5 word554 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3867 Y6 word606 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3868 GND word951 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3869 Y7 word892 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3870 Y1 word152 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3871 GND word371 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3872 Y7 word210 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3873 Y1 word640 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3874 Y0 word658 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3875 Y2 word936 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3876 GND word995 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X3877 GND word743 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3878 Y7 word146 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3879 Y2 word834 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X3880 GND word883 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3881 GND word711 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3882 GND word939 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X3883 GND word251 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3884 Y5 word370 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3885 Y1 word520 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3886 GND word579 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3887 Y5 word700 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3888 Y5 word148 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3889 GND word307 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X3890 GND word875 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3891 GND word205 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3892 Y1 word298 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3893 Y1 word628 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3894 Y5 word636 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3895 GND word137 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3896 GND word141 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3897 GND word763 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3898 Y1 word684 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3899 Y2 word412 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X3900 Y5 word682 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3901 Y2 word678 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3902 GND word187 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3903 GND word735 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3904 GND word159 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3905 GND word453 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3906 Y3 word604 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3907 GND word663 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3908 Y0 word744 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3909 Y2 word558 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3910 Y1 word776 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3911 Y4 word166 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3912 Y0 word1010 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3913 GND word157 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3914 Y0 word316 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3915 GND word471 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3916 GND word881 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X3917 Y4 word722 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3918 Y0 word150 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3919 GND word271 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3920 GND word305 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3921 Y5 word874 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3922 Y6 word246 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3923 GND word421 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3924 GND word203 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3925 Y3 word262 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X3926 GND word357 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3927 Y0 word992 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X3928 GND word255 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3929 Y7 word916 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3930 GND word857 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3931 GND word827 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3932 Y0 word196 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3933 Y6 word410 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3934 Y3 word528 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3935 Y4 word534 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3936 GND word755 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3937 GND word525 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3938 GND word863 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3939 GND word253 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3940 GND word303 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X3941 Y0 word462 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3942 GND word617 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3943 Y1 word968 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3944 GND word237 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3945 Y0 word296 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3946 GND word961 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X3947 Y6 word392 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3948 GND word417 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3949 GND word451 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3950 GND word575 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3951 Y4 word634 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3952 GND word737 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3953 Y7 word216 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3954 Y2 word904 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3955 GND word869 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3956 GND word503 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X3957 Y5 word174 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3958 Y4 word192 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3959 GND word973 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3960 GND word781 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3961 Y0 word342 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X3962 GND word321 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3963 Y3 word950 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3964 GND word1009 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3965 Y7 word842 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3966 Y6 word974 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3967 GND word915 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3968 GND word279 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3969 Y0 word608 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X3970 GND word945 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.2193 ps=1.88 w=0.51 l=0.17
X3971 Y3 word784 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X3972 GND word155 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3973 GND word749 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3974 GND word207 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3975 GND word215 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3976 Y1 word424 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3977 Y2 word152 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3978 GND word545 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3979 GND word991 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X3980 Y2 word720 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3981 GND word695 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X3982 GND word143 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3983 Y7 word362 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3984 Y2 word640 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3985 GND word889 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3986 Y3 word830 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X3987 GND word201 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X3988 Y5 word320 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X3989 GND word927 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X3990 Y2 word986 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4635 ps=3.36 w=0.51 l=0.17
X3991 Y1 word470 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X3992 GND word689 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X3993 Y1 word248 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3994 Y7 word408 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3995 Y7 word242 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3996 Y2 word520 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X3997 Y0 word814 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4635 ps=3.36 w=0.51 l=0.17
X3998 Y5 word632 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X3999 GND word691 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4000 GND word137 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4001 Y5 word568 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4002 Y3 word224 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4003 Y3 word554 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4004 Y6 word316 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4005 GND word885 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4006 GND word673 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X4007 GND word897 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4008 Y6 word150 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4009 Y0 word266 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X4010 Y4 word604 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4011 Y4 word894 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4012 Y7 word766 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4013 GND word933 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X4014 GND word357 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4015 GND word255 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X4016 Y5 word824 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4017 GND word765 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4018 Y6 word196 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4019 GND word379 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4020 Y1 word708 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X4021 GND word157 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4022 GND word307 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X4023 Y0 word366 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X4024 Y3 word700 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X4025 Y3 word148 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4026 GND word205 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4027 Y6 word462 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4028 Y7 word866 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4029 Y4 word484 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4030 Y3 word636 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X4031 GND word475 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X4032 GND word813 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X4033 GND word141 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4034 GND word203 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4035 GND word237 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4036 Y6 word296 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4037 Y5 word806 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4038 Y0 word412 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X4039 Y0 word570 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X4040 Y7 word912 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4041 Y6 word714 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4042 Y3 word682 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4043 Y4 word818 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4044 GND word187 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4045 GND word911 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4046 Y7 word848 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4047 Y0 word678 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X4048 GND word921 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4049 GND word795 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4050 Y7 word166 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4051 GND word819 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4052 Y6 word760 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4053 GND word285 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4054 GND word303 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4055 GND word453 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X4056 Y7 word654 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4057 Y1 word274 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4058 Y6 word608 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4059 GND word953 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4060 Y4 word630 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4061 Y3 word900 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4062 Y5 word390 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4063 GND word429 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4064 Y1 word540 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X4065 Y0 word558 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X4066 GND word895 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4067 Y6 word860 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4068 Y2 word836 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X4069 Y3 word734 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4070 GND word165 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4071 Y1 word374 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4072 GND word941 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X4073 GND word253 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4074 Y2 word590 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4075 GND word965 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4076 Y6 word906 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4077 Y5 word372 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4078 GND word431 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X4079 GND word149 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4080 GND word211 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4081 Y5 word702 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4082 GND word207 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4083 Y1 word420 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4084 Y1 word198 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4085 Y2 word424 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X4086 Y5 word638 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4087 Y1 word356 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4088 GND word417 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4089 GND word695 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4090 GND word143 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4091 GND word353 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X4092 Y2 word982 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4093 Y7 word192 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4094 GND word683 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4095 GND word311 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4096 Y2 word918 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X4097 Y0 word764 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X4098 Y7 word680 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4099 Y2 word248 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4100 GND word971 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X4101 Y1 word668 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X4102 Y4 word964 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4103 Y3 word174 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4104 GND word623 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4105 GND word805 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.2193 ps=1.88 w=0.51 l=0.17
X4106 Y0 word746 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X4107 Y3 word440 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X4108 GND word279 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X4109 Y0 word1012 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X4110 Y4 word224 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4111 GND word215 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4112 Y0 word152 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4113 GND word307 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4114 Y6 word366 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4115 GND word939 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.2193 ps=1.88 w=0.51 l=0.17
X4116 Y5 word876 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4117 GND word205 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4118 Y0 word640 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X4119 GND word329 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X4120 Y3 word320 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X4121 Y4 word888 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4122 GND word141 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4123 GND word257 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X4124 Y6 word412 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4125 GND word951 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.2193 ps=1.88 w=0.51 l=0.17
X4126 GND word595 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4127 Y4 word944 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X4128 GND word757 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4129 GND word527 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4130 Y3 word586 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4131 GND word917 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X4132 GND word763 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X4133 GND word187 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4134 Y5 word756 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4135 Y0 word520 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X4136 Y4 word700 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4137 Y4 word148 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4138 Y0 word298 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2914 ps=1.87 w=0.51 l=0.17
X4139 GND word453 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4140 Y4 word636 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4141 GND word963 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4142 GND word137 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4143 Y0 word628 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X4144 VDD GND Y4 VDD sky130_fd_pr__pfet_01v8 ad=0.1836 pd=1.74 as=0.1836 ps=1.74 w=0.51 l=0.17
X4145 GND word871 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4146 Y3 word804 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X4147 GND word745 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X4148 Y0 word684 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.40905 ps=2.7 w=0.51 l=0.17
X4149 GND word235 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4150 GND word403 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4371 pd=2.81 as=0.1377 ps=1.05 w=0.51 l=0.17
X4151 GND word903 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4152 GND word705 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X4153 Y6 word976 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4154 GND word909 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4155 GND word219 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4156 Y1 word160 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4157 GND word281 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2931 pd=1.88 as=0.1377 ps=1.05 w=0.51 l=0.17
X4158 Y5 word340 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
X4159 GND word379 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4160 Y1 word490 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4161 GND word947 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X4162 Y3 word786 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4163 GND word157 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4164 GND word217 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4165 GND word751 Y6 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4166 Y1 word426 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4167 GND word547 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4168 GND word645 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4169 Y1 word324 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4170 GND word891 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4171 GND word203 Y7 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4172 GND word381 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4173 GND word531 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X4174 Y2 word988 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.3101 ps=1.945 w=0.51 l=0.17
X4175 Y5 word156 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4176 GND word315 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X4177 Y1 word306 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4178 Y5 word486 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4179 GND word873 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4180 GND word149 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4181 GND word581 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X4182 Y0 word816 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2914 ps=1.87 w=0.51 l=0.17
X4183 Y2 word420 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.2598 ps=1.79 w=0.51 l=0.17
X4184 Y1 word572 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X4185 GND word809 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4186 GND word693 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4187 Y2 word198 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4188 Y2 word356 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X4189 Y2 word686 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4190 GND word285 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X4191 Y4 word914 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4192 GND word857 Y0 GND sky130_fd_pr__nfet_01v8 ad=0.4116 pd=2.71 as=0.1377 ps=1.05 w=0.51 l=0.17
X4193 GND word461 Y2 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.2193 ps=1.88 w=0.51 l=0.17
X4194 Y1 word950 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X4195 Y4 word850 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4196 Y1 word728 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.40905 ps=2.7 w=0.51 l=0.17
X4197 Y6 word152 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4198 Y0 word962 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.4116 ps=2.71 w=0.51 l=0.17
X4199 Y1 word784 GND GND sky130_fd_pr__nfet_01v8 ad=0.2244 pd=1.9 as=0.43965 ps=2.82 w=0.51 l=0.17
X4200 Y4 word174 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.3101 ps=1.945 w=0.51 l=0.17
X4201 Y6 word640 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.4116 ps=2.71 w=0.51 l=0.17
X4202 GND word165 Y3 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.1377 ps=1.05 w=0.51 l=0.17
X4203 GND word833 Y1 GND sky130_fd_pr__nfet_01v8 ad=0.41415 pd=2.72 as=0.1377 ps=1.05 w=0.51 l=0.17
X4204 Y0 word796 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X4205 GND word733 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.2598 pd=1.79 as=0.1377 ps=1.05 w=0.51 l=0.17
X4206 Y5 word826 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.43965 ps=2.82 w=0.51 l=0.17
X4207 GND word789 Y4 GND sky130_fd_pr__nfet_01v8 ad=0.4686 pd=3.38 as=0.1377 ps=1.05 w=0.51 l=0.17
X4208 GND word767 Y5 GND sky130_fd_pr__nfet_01v8 ad=0.3101 pd=1.945 as=0.2193 ps=1.88 w=0.51 l=0.17
X4209 Y4 word730 GND GND sky130_fd_pr__nfet_01v8 ad=0.1377 pd=1.05 as=0.2598 ps=1.79 w=0.51 l=0.17
.ends

.subckt mux2 I1 I0 S0 VDD GND Y ~S0
X0 GND I0 a_72_226# GND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.89 as=0.18 ps=1.72 w=0.5 l=0.15
X1 a_72_226# S0 GND GND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.89 as=0.0975 ps=0.89 w=0.5 l=0.15
X2 Y ~S0 a_72_226# GND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.89 as=0.0975 ps=0.89 w=0.5 l=0.15
X3 a_174_630# I0 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X4 Y S0 a_174_630# VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X5 a_72_226# I1 Y GND sky130_fd_pr__nfet_01v8 ad=0.18 pd=1.72 as=0.0975 ps=0.89 w=0.5 l=0.15
X6 a_390_630# ~S0 Y VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7 VDD I1 a_390_630# VDD sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.72 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt mux4 I1 I2 I3 S0 ~S0 S1 ~S1 Y VDD I0 GND
Xmux2_0 I1 I0 S0 VDD GND mux2_0/Y ~S0 mux2
Xmux2_1 I3 I2 S0 VDD GND mux2_1/Y ~S0 mux2
Xmux2_2 mux2_1/Y mux2_0/Y S1 VDD GND Y ~S1 mux2
.ends

.subckt inv VDD GND A Y
X0 Y A GND GND sky130_fd_pr__nfet_01v8 ad=0.18 pd=1.72 as=0.18 ps=1.72 w=0.5 l=0.15
X1 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.72 as=0.36 ps=2.72 w=1 l=0.15
.ends

.subckt nand VDD GND A Y B
X0 a_174_130# B GND GND sky130_fd_pr__nfet_01v8 ad=0.0525 pd=0.71 as=0.18 ps=1.72 w=0.5 l=0.15
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 VDD A Y VDD sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.72 as=0.195 ps=1.39 w=1 l=0.15
X3 Y A a_174_130# GND sky130_fd_pr__nfet_01v8 ad=0.18 pd=1.72 as=0.0525 ps=0.71 w=0.5 l=0.15
.ends

.subckt dff D ~CLK CLK ~Q Q VDD GND
X0 ~Q Q VDD VDD sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.72 as=0.195 ps=1.39 w=1 l=0.15
X1 a_174_130# ~CLK D GND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.89 as=0.18 ps=1.72 w=0.5 l=0.15
X2 VDD a_174_130# a_422_130# VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X3 a_282_130# CLK a_174_130# GND sky130_fd_pr__nfet_01v8 ad=0.18 pd=1.72 as=0.0975 ps=0.89 w=0.5 l=0.15
X4 a_282_130# a_422_130# GND GND sky130_fd_pr__nfet_01v8 ad=0.18 pd=1.72 as=0.0975 ps=0.89 w=0.5 l=0.15
X5 a_174_130# CLK D VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X6 a_282_130# ~CLK a_174_130# VDD sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.72 as=0.195 ps=1.39 w=1 l=0.15
X7 a_282_130# a_422_130# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.72 as=0.195 ps=1.39 w=1 l=0.15
X8 a_906_130# CLK a_422_130# GND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.89 as=0.18 ps=1.72 w=0.5 l=0.15
X9 ~Q ~CLK a_906_130# GND sky130_fd_pr__nfet_01v8 ad=0.18 pd=1.72 as=0.0975 ps=0.89 w=0.5 l=0.15
X10 GND a_906_130# Q GND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.89 as=0.18 ps=1.72 w=0.5 l=0.15
X11 a_906_130# ~CLK a_422_130# VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X12 ~Q Q GND GND sky130_fd_pr__nfet_01v8 ad=0.18 pd=1.72 as=0.0975 ps=0.89 w=0.5 l=0.15
X13 GND a_174_130# a_422_130# GND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.89 as=0.18 ps=1.72 w=0.5 l=0.15
X14 ~Q CLK a_906_130# VDD sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.72 as=0.195 ps=1.39 w=1 l=0.15
X15 VDD a_906_130# Q VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
.ends

.subckt xor VDD GND Y A ~B ~A B
X0 Y ~A a_300_226# GND sky130_fd_pr__nfet_01v8 ad=0.095 pd=0.88 as=0.0525 ps=0.71 w=0.5 l=0.15
X1 GND A a_90_226# GND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.89 as=0.18 ps=1.72 w=0.5 l=0.15
X2 VDD B a_390_630# VDD sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.72 as=0.105 ps=1.21 w=1 l=0.15
X3 a_300_226# ~B GND GND sky130_fd_pr__nfet_01v8 ad=0.0525 pd=0.71 as=0.0975 ps=0.89 w=0.5 l=0.15
X4 Y ~B a_210_630# VDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X5 a_390_630# ~A Y VDD sky130_fd_pr__pfet_01v8 ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X6 a_210_630# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.105 pd=1.21 as=0.36 ps=2.72 w=1 l=0.15
X7 a_90_226# B Y GND sky130_fd_pr__nfet_01v8 ad=0.18 pd=1.72 as=0.095 ps=0.88 w=0.5 l=0.15
.ends

.subckt tff T CLK ~CLK Q ~Q xor_0/GND VDD
Xdff_0 xor_0/Y ~CLK CLK ~Q Q VDD xor_0/GND dff
Xxor_0 VDD xor_0/GND xor_0/Y T ~Q inv_0/Y Q xor
Xinv_0 VDD xor_0/GND T inv_0/Y inv
.ends

.subckt counter_8 CLK Q0 Q2 Q3 Q4 Q5 Q6 Q7 GND Q1 VDD
Xnand_3 VDD GND tff_5/T inv_0/A Q6 nand
Xnand_4 VDD GND tff_6/T inv_5/A Q5 nand
Xnand_5 VDD GND tff_7/T inv_6/A Q4 nand
Xnand_6 VDD GND tff_4/T inv_7/A Q3 nand
Xtff_0 tff_0/T CLK inv_1/Y Q2 tff_0/~Q GND VDD tff
Xtff_1 VDD CLK inv_1/Y Q0 tff_1/~Q GND VDD tff
Xtff_2 tff_2/T CLK inv_1/Y Q1 tff_2/~Q GND VDD tff
Xtff_3 tff_3/T CLK inv_1/Y Q7 tff_3/~Q GND VDD tff
Xtff_4 tff_4/T CLK inv_1/Y Q3 tff_4/~Q GND VDD tff
Xtff_5 tff_5/T CLK inv_1/Y Q6 tff_5/~Q GND VDD tff
Xtff_6 tff_6/T CLK inv_1/Y Q5 tff_6/~Q GND VDD tff
Xtff_7 tff_7/T CLK inv_1/Y Q4 tff_7/~Q GND VDD tff
Xinv_0 VDD GND inv_0/A tff_3/T inv
Xinv_1 VDD GND CLK inv_1/Y inv
Xinv_2 VDD GND inv_2/A tff_2/T inv
Xinv_3 VDD GND inv_3/A tff_0/T inv
Xinv_4 VDD GND inv_4/A tff_4/T inv
Xinv_5 VDD GND inv_5/A tff_5/T inv
Xinv_6 VDD GND inv_6/A tff_6/T inv
Xinv_7 VDD GND inv_7/A tff_7/T inv
Xnand_0 VDD GND tff_0/T inv_4/A Q2 nand
Xnand_1 VDD GND VDD inv_2/A Q0 nand
Xnand_2 VDD GND tff_2/T inv_3/A Q1 nand
.ends

.subckt decoder_8 A0 A1 A2 A3 A4 A5 A6 word0 word1 word2 word3 word4 word5 word6 word7
+ word8 word9 word10 word11 word12 word13 word14 word15 word16 word17 word18 word19
+ word20 word21 word22 word23 word24 word25 word26 word27 word28 word29 word30 word31
+ word32 word33 word34 word35 word36 word37 word38 word39 word40 word41 word42 word43
+ word44 word45 word46 word47 word48 word49 word50 word51 word52 word53 word54 word55
+ word56 word57 word58 word59 word60 word61 word62 word63 word64 word65 word66 word67
+ word68 word69 word70 word71 word72 word73 word74 word75 word76 word77 word78 word79
+ word80 word81 word82 word83 word84 word85 word86 word87 word88 word89 word90 word91
+ word92 word93 word94 word95 word96 word97 word98 word99 word100 word101 word102
+ word103 word104 word105 word106 word107 word108 word109 word110 word111 word112
+ word113 word114 word115 word116 word117 word118 word119 word120 word121 word122
+ word123 word124 word125 word126 word127 word128 word129 word130 word131 word132
+ word133 word134 word135 word136 word137 word138 word139 word140 word141 word142
+ word143 word144 word145 word146 word147 word148 word149 word150 word151 word152
+ word153 word154 word155 word156 word157 word158 word159 word160 word161 word162
+ word163 word164 word165 word166 word167 word168 word169 word170 word171 word172
+ word173 word174 word175 word176 word177 word178 word179 word180 word181 word182
+ word183 word184 word185 word186 word187 word188 word189 word190 word191 word192
+ word193 word194 word195 word196 word197 word198 word199 word200 word201 word202
+ word203 word204 word205 word206 word207 word208 word209 word210 word211 word212
+ word213 word214 word215 word216 word217 word218 word219 word220 word221 word222
+ word223 word224 word225 word226 word227 word228 word229 word230 word231 word232
+ word233 word234 word235 word236 word237 word238 word239 word240 word241 word242
+ word243 word244 word245 word246 word247 word248 word249 word250 word251 word252
+ word253 word254 word255 word256 word257 word258 word259 word260 word261 word262
+ word263 word264 word265 word266 word267 word268 word269 word270 word271 word272
+ word273 word274 word275 word276 word277 word278 word279 word280 word281 word282
+ word283 word284 word285 word286 word287 word288 word289 word290 word291 word292
+ word293 word294 word295 word296 word297 word298 word299 word300 word301 word302
+ word303 word304 word305 word306 word307 word308 word309 word310 word311 word312
+ word313 word314 word315 word316 word317 word318 word319 word320 word321 word322
+ word323 word324 word325 word326 word327 word328 word329 word330 word331 word332
+ word333 word334 word335 word336 word337 word338 word339 word340 word341 word342
+ word343 word344 word345 word346 word347 word348 word349 word350 word351 word352
+ word353 word354 word355 word356 word357 word358 word359 word360 word361 word362
+ word363 word364 word365 word366 word367 word368 word369 word370 word371 word372
+ word373 word374 word375 word376 word377 word378 word379 word380 word381 word382
+ word383 word384 word385 word386 word387 word388 word389 word390 word391 word392
+ word393 word394 word395 word396 word397 word398 word399 word400 word401 word402
+ word403 word404 word405 word406 word407 word408 word409 word410 word411 word412
+ word413 word414 word415 word416 word417 word418 word419 word420 word421 word422
+ word423 word424 word425 word426 word427 word428 word429 word430 word431 word432
+ word433 word434 word435 word436 word437 word438 word439 word440 word441 word442
+ word443 word444 word445 word446 word447 word448 word449 word450 word451 word452
+ word453 word454 word455 word456 word457 word458 word459 word460 word461 word462
+ word463 word464 word465 word466 word467 word468 word469 word470 word471 word472
+ word473 word474 word475 word476 word477 word478 word479 word480 word481 word482
+ word483 word484 word485 word486 word487 word488 word489 word490 word491 word492
+ word493 word494 word495 word496 word497 word498 word499 word500 word501 word502
+ word503 word504 word505 word506 word507 word508 word509 word510 word511 word512
+ word513 word514 word515 word516 word517 word518 word519 word520 word521 word522
+ word523 word524 word525 word526 word527 word528 word529 word530 word531 word532
+ word533 word534 word535 word536 word537 word538 word539 word540 word541 word542
+ word543 word544 word545 word546 word547 word548 word549 word550 word551 word552
+ word553 word554 word555 word556 word557 word558 word559 word560 word561 word562
+ word563 word564 word565 word566 word567 word568 word569 word570 word571 word572
+ word573 word574 word575 word576 word577 word578 word579 word580 word581 word582
+ word583 word584 word585 word586 word587 word588 word589 word590 word591 word592
+ word593 word594 word595 word596 word597 word598 word599 word600 word601 word602
+ word603 word604 word605 word606 word607 word608 word609 word610 word611 word612
+ word613 word614 word615 word616 word617 word618 word619 word620 word621 word622
+ word623 word624 word625 word626 word627 word628 word629 word630 word631 word632
+ word633 word634 word635 word636 word637 word638 word639 word640 word641 word642
+ word643 word644 word645 word646 word647 word648 word649 word650 word651 word652
+ word653 word654 word655 word656 word657 word658 word659 word660 word661 word662
+ word663 word664 word665 word666 word667 word668 word669 word670 word671 word672
+ word673 word674 word675 word676 word677 word678 word679 word680 word681 word682
+ word683 word684 word685 word686 word687 word688 word689 word690 word691 word692
+ word693 word694 word695 word696 word697 word698 word699 word700 word701 word702
+ word703 word704 word705 word706 word707 word708 word709 word710 word711 word712
+ word713 word714 word715 word716 word717 word718 word719 word720 word721 word722
+ word723 word724 word725 word726 word727 word728 word729 word730 word731 word732
+ word733 word734 word735 word736 word737 word738 word739 word740 word741 word742
+ word743 word744 word745 word746 word747 word748 word749 word750 word751 word752
+ word753 word754 word755 word756 word757 word758 word759 word760 word761 word762
+ word763 word764 word765 word766 word767 word768 word769 word770 word771 word772
+ word773 word774 word775 word776 word777 word778 word779 word780 word781 word782
+ word783 word784 word785 word786 word787 word788 word789 word790 word791 word792
+ word793 word794 word795 word796 word797 word798 word799 word800 word801 word802
+ word803 word804 word805 word806 word807 word808 word809 word810 word811 word812
+ word813 word814 word815 word816 word817 word818 word819 word820 word821 word822
+ word823 word824 word825 word826 word827 word828 word829 word830 word831 word832
+ word833 word834 word835 word836 word837 word838 word839 word840 word841 word842
+ word843 word844 word845 word846 word847 word848 word849 word850 word851 word852
+ word853 word854 word855 word856 word857 word858 word859 word860 word861 word862
+ word863 word864 word865 word866 word867 word868 word869 word870 word871 word872
+ word873 word874 word875 word876 word877 word878 word879 word880 word881 word882
+ word883 word884 word885 word886 word887 word888 word889 word890 word891 word892
+ word893 word894 word895 word896 word897 word898 word899 word900 word901 word902
+ word903 word904 word905 word906 word907 word908 word909 word910 word911 word912
+ word913 word914 word915 word916 word917 word918 word919 word920 word921 word922
+ word923 word924 word925 word926 word927 word928 word929 word930 word931 word932
+ word933 word934 word935 word936 word937 word938 word939 word940 word941 word942
+ word943 word944 word945 word946 word947 word948 word949 word950 word951 word952
+ word953 word954 word955 word956 word957 word958 word959 word960 word961 word962
+ word963 word964 word965 word966 word967 word968 word969 word970 word971 word972
+ word973 word974 word975 word976 word977 word978 word979 word980 word981 word982
+ word983 word984 word985 word986 word987 word988 word989 word990 word991 word992
+ word993 word994 word995 word996 word997 word998 word999 word1000 word1001 word1002
+ word1003 word1004 word1005 word1006 word1007 word1008 word1009 word1010 word1011
+ word1012 word1013 word1014 word1015 word1016 word1017 word1018 word1019 word1020
+ word1021 word1022 word1023 VDD GND A7 A8 A9
X0 a_578_n94630# a_528_n66# a_446_n94630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1 word703 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2 word357 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3 word694 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4 a_578_n33286# a_528_n66# a_446_n33286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5 a_842_n104996# a_792_n66# a_578_n104996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6 word9 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7 word260 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8 word974 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9 a_1766_n143904# A3 a_1370_n143904# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10 GND A3 word166 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11 a_1106_n88098# a_1056_n66# a_842_n88098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12 a_2294_n13832# A1 a_2030_n13832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13 a_314_n116782# a_264_n66# a_50_n116782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14 GND A6 word538 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15 word999 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16 word91 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17 word940 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18 a_314_n53450# a_264_n66# a_182_n53450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19 a_1634_n103718# a_1584_n66# a_1370_n103718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20 a_974_n117634# A6 a_710_n117634# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X21 word316 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X22 GND A0 word540 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X23 word836 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X24 word465 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X25 a_182_n23488# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X26 a_842_n89376# a_792_n66# a_710_n89376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X27 a_578_n71058# a_528_n66# a_314_n71058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X28 GND A3 word274 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X29 a_1898_n53166# a_1848_n66# a_1766_n53166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X30 a_842_n142768# a_792_n66# a_578_n142768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X31 word819 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X32 a_578_n62680# a_528_n66# a_314_n62680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X33 word469 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X34 word528 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X35 word764 A0 a_2294_n108688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X36 GND A3 word432 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X37 word217 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X38 word486 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X39 a_1502_n74892# A4 a_1238_n74892# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X40 GND A2 word880 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X41 a_1766_n111954# A3 a_1370_n111954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X42 a_710_n17808# A7 a_446_n17808# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X43 word749 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X44 a_1238_n38114# A5 a_974_n38114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X45 word530 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X46 a_1238_n29736# A5 a_842_n29736# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X47 a_2294_n28742# A1 a_2030_n28742# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X48 a_1634_n77306# a_1584_n66# a_1370_n77306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X49 a_2162_n21642# a_2112_n66# a_1898_n21642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X50 a_182_n61260# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X51 a_314_n68360# a_264_n66# a_182_n68360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X52 word137 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X53 GND A3 word210 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X54 a_1634_n127006# a_1584_n66# a_1370_n127006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X55 a_314_n123030# a_264_n66# a_50_n123030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X56 a_1106_n126438# a_1056_n66# a_842_n126438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X57 word363 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X58 word422 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X59 a_1898_n82560# a_1848_n66# a_1766_n82560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X60 GND A5 word89 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X61 GND A5 word148 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X62 a_1238_n20648# A5 a_974_n20648# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X63 word356 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X64 a_182_n38398# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X65 word266 A0 a_2162_n37972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X66 word1015 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X67 GND A9 word141 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X68 word505 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X69 GND A9 word82 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X70 word202 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X71 a_1238_n67508# A5 a_842_n67508# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X72 a_1898_n68076# a_1848_n66# a_1634_n68076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X73 word686 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X74 word73 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X75 GND A9 word412 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X76 GND A1 word736 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X77 a_1766_n135242# A3 a_1370_n135242# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X78 a_1634_n45356# a_1584_n66# a_1370_n45356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X79 word403 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X80 GND A0 word640 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X81 word877 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X82 word628 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X83 GND A0 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X84 word527 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X85 word532 A0 a_2294_n75744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X86 word689 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X87 word345 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X88 a_2030_n135810# A2 a_1634_n135810# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X89 word941 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X90 GND A0 word28 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X91 word38 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X92 a_2030_n14116# A2 a_1766_n14116# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X93 a_1898_n97470# a_1848_n66# a_1634_n97470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X94 word790 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X95 GND A5 word194 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X96 a_4084_164# A4 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X97 word470 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X98 GND A9 word246 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X99 GND A9 word187 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X100 a_1634_n74750# a_1584_n66# a_1502_n74750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X101 word564 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X102 a_1634_n83128# a_1584_n66# a_1502_n83128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X103 a_2030_n83412# A2 a_1634_n83412# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X104 a_1766_n103292# A3 a_1370_n103292# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X105 a_2030_n143762# A2 a_1766_n143762# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X106 word310 A0 a_2162_n44220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X107 GND A8 word86 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X108 a_2162_n74324# a_2112_n66# a_2030_n74324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X109 word996 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X110 a_1106_n132260# a_1056_n66# a_974_n132260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X111 word711 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X112 a_1634_n124450# a_1584_n66# a_1502_n124450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X113 GND A1 word841 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X114 a_2162_n65946# a_2112_n66# a_1898_n65946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X115 a_446_n105422# A8 a_50_n105422# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X116 word239 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X117 a_710_n78442# A7 a_446_n78442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X118 a_974_n129988# A6 a_578_n129988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X119 word180 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X120 a_1502_n96050# A4 a_1106_n96050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X121 word982 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X122 a_2030_n43510# A2 a_1766_n43510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X123 word366 A0 a_2162_n52172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X124 a_578_n105706# a_528_n66# a_446_n105706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X125 a_2030_n103860# A2 a_1634_n103860# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X126 word302 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X127 GND A5 word460 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X128 word464 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X129 a_1238_n73330# A5 a_974_n73330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X130 word696 A0 a_2294_n99032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X131 word715 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X132 GND A9 word453 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X133 GND A3 word519 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X134 GND A3 word578 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X135 GND A6 word916 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X136 a_1766_n141064# A3 a_1502_n141064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X137 a_2030_n29026# A2 a_1634_n29026# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X138 a_2294_n63958# A1 a_2030_n63958# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X139 a_2294_n72336# A1 a_1898_n72336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X140 GND A3 word722 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X141 a_1766_n132686# A3 a_1502_n132686# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X142 GND A1 word777 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X143 a_710_n38540# A7 a_314_n38540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X144 word245 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X145 word895 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X146 word760 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X147 word781 a_2376_n66# a_2294_n111102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X148 a_1634_n42800# a_1584_n66# a_1502_n42800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X149 a_2030_n51462# A2 a_1634_n51462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X150 word385 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X151 GND A5 word516 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X152 a_2162_n105138# a_2112_n66# a_2030_n105138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X153 word669 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X154 a_1898_n132970# a_1848_n66# a_1766_n132970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X155 a_446_n15820# A8 a_182_n15820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X156 a_2030_n89944# A2 a_1634_n89944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X157 a_710_n113942# A7 a_314_n113942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X158 a_2030_n98322# A2 a_1766_n98322# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X159 a_2162_n33996# a_2112_n66# a_1898_n33996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X160 a_710_n46492# A7 a_314_n46492# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X161 a_1502_n64100# A4 a_1238_n64100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X162 GND A8 word191 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X163 a_2162_n89234# a_2112_n66# a_2030_n89234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X164 word757 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X165 word765 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X166 GND A8 word132 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X167 a_1766_n75602# A3 a_1370_n75602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X168 a_2030_n11560# A2 a_1766_n11560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X169 word502 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X170 a_446_n23772# A8 a_182_n23772# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X171 GND A6 word61 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X172 GND A7 word818 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X173 a_1106_n5738# a_1056_n66# a_974_n5738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X174 GND A2 word193 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X175 a_2030_n58420# A2 a_1634_n58420# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X176 GND A9 word228 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X177 a_2030_n118770# A2 a_1766_n118770# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X178 word821 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X179 a_2030_n80856# A2 a_1634_n80856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X180 GND A5 word133 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X181 word219 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X182 a_2162_n80146# a_2112_n66# a_2030_n80146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X183 a_2294_n87246# A1 a_1898_n87246# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X184 GND A2 word681 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X185 GND A3 word886 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X186 a_2294_n100310# A1 a_2030_n100310# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X187 GND A9 word126 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X188 a_2030_n66372# A2 a_1766_n66372# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X189 word350 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X190 a_710_n84264# A7 a_446_n84264# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X191 a_446_n102866# A8 a_50_n102866# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X192 word549 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X193 word827 a_2376_n66# a_2162_n117634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X194 VDD A3 a_1584_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X195 a_710_n75886# A7 a_446_n75886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X196 word1023 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X197 word190 A0 a_2162_n27180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X198 a_2162_n142484# a_2112_n66# a_2030_n142484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X199 word791 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X200 word829 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X201 a_974_n6022# A6 a_710_n6022# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X202 a_2162_n57284# a_2112_n66# a_2030_n57284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X203 GND A1 word60 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X204 a_1766_n43652# A3 a_1370_n43652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X205 word119 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X206 word678 A0 a_2162_n96476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X207 GND A9 word494 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X208 GND A5 word793 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X209 a_1106_n33002# a_1056_n66# a_842_n33002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X210 GND A9 word435 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X211 a_1106_n24624# a_1056_n66# a_974_n24624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X212 GND A8 word15 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X213 word614 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X214 a_2030_n26470# A2 a_1634_n26470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X215 GND A5 word340 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X216 word303 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X217 a_1238_n56290# A5 a_974_n56290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X218 word1017 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X219 GND A9 word333 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X220 a_446_n30020# A8 a_182_n30020# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X221 a_1766_n12128# A3 a_1370_n12128# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X222 a_2294_n55296# A1 a_1898_n55296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X223 GND A2 word456 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X224 a_2030_n95766# A2 a_1766_n95766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X225 GND A0 word986 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X226 word865 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X227 GND A8 word173 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X228 GND A8 word232 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X229 GND A7 word517 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X230 GND A8 word734 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X231 word65 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X232 a_1238_n129562# A5 a_974_n129562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X233 a_2294_n910# A1 a_1898_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X234 word81 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X235 a_446_n90938# A8 a_50_n90938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X236 GND A7 word34 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X237 a_446_n626# A8 a_182_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X238 GND A2 word234 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X239 GND A7 word800 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X240 GND A7 word859 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X241 GND A9 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X242 a_1370_n129846# a_1320_n66# a_1238_n129846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X243 GND A0 word766 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X244 a_446_n5312# A8 a_182_n5312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X245 a_446_n76454# A8 a_50_n76454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X246 word510 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X247 GND A5 word898 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X248 a_1502_n138508# A4 a_1238_n138508# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X249 word78 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X250 a_974_n23914# A6 a_578_n23914# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X251 word851 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X252 word450 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X253 word792 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X254 GND A3 word868 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X255 GND A1 word864 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X256 a_1238_n120474# A5 a_842_n120474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X257 a_2030_n72194# A2 a_1634_n72194# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X258 a_710_n90086# A7 a_446_n90086# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X259 a_1370_n80004# a_1320_n66# a_1106_n80004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X260 word349 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X261 word408 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X262 a_1370_n71626# a_1320_n66# a_1106_n71626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X263 word279 a_2376_n66# a_2162_n39818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X264 GND A7 word351 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X265 GND A2 word561 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X266 a_1370_n120758# a_1320_n66# a_1238_n120758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X267 a_1898_n1904# a_1848_n66# a_1634_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X268 a_1766_n18660# A3 a_1502_n18660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X269 GND A7 word292 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X270 a_974_n3466# A6 a_710_n3466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X271 GND A1 word432 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X272 GND A9 word49 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X273 a_1370_n48764# a_1320_n66# a_1238_n48764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X274 a_1370_n57142# a_1320_n66# a_1238_n57142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X275 GND A7 word622 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X276 a_1766_n96334# A3 a_1502_n96334# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X277 GND A5 word29 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X278 word186 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X279 word926 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X280 GND A5 word732 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X281 word285 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X282 GND A2 word339 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X283 a_1106_n68928# a_1056_n66# a_842_n68928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X284 GND A4 word770 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X285 word215 a_2376_n66# a_2162_n30730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X286 GND A7 word70 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X287 GND A2 word280 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X288 a_1502_n106558# A4 a_1106_n106558# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X289 word64 A0 a_2294_n9288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X290 GND A2 word497 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X291 GND A4 word928 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X292 a_1370_n17240# a_1320_n66# a_1106_n17240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X293 GND A0 word810 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X294 GND A5 word26 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X295 word113 a_2376_n66# a_2294_n16246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X296 a_842_n31724# a_792_n66# a_578_n31724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X297 word181 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X298 a_974_n38824# A6 a_710_n38824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X299 GND A8 word214 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X300 a_2294_n99600# A1 a_1898_n99600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X301 a_1766_n2614# A3 a_1370_n2614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X302 a_2162_n7868# a_2112_n66# a_1898_n7868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X303 a_2162_n92500# a_2112_n66# a_2030_n92500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X304 word897 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X305 word973 a_2376_n66# a_2294_n138366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X306 GND A1 word969 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X307 GND A3 word914 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X308 word762 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X309 GND A8 word544 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X310 a_1370_n25192# a_1320_n66# a_1106_n25192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X311 word671 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X312 word743 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X313 a_1370_n144046# a_1320_n66# a_1106_n144046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X314 word975 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X315 GND A0 word866 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X316 word601 a_2376_n66# a_2294_n85542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X317 a_1370_n135668# a_1320_n66# a_1106_n135668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X318 a_578_n132260# a_528_n66# a_314_n132260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X319 a_50_n134532# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X320 a_446_n82276# A8 a_50_n82276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X321 GND A1 word537 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X322 a_446_n2756# A8 a_182_n2756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X323 a_446_n73898# A8 a_50_n73898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X324 a_1766_n64384# A3 a_1502_n64384# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X325 a_1106_n45356# a_1056_n66# a_974_n45356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X326 GND A2 word114 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X327 GND A6 word296 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X328 GND A3 word850 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X329 a_710_n1052# A7 a_446_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X330 a_50_n90512# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X331 GND A5 word837 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X332 word379 a_2376_n66# a_2162_n54018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X333 a_50_n103008# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X334 a_2294_n4744# A1 a_2030_n4744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X335 GND A0 word298 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X336 GND A2 word602 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X337 a_710_n118060# A7 a_314_n118060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X338 GND A2 word801 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X339 GND A4 word291 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X340 a_1370_n54586# a_1320_n66# a_1106_n54586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X341 a_842_n46634# a_792_n66# a_710_n46634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X342 GND A7 word604 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X343 word862 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X344 word809 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X345 a_1238_n1904# A5 a_974_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X346 GND A0 word196 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X347 a_1766_n93778# A3 a_1370_n93778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X348 a_1370_n112096# a_1320_n66# a_1238_n112096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X349 word750 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X350 a_182_n27606# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X351 a_50_n102582# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X352 a_314_n111812# a_264_n66# a_50_n111812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X353 GND A6 word562 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X354 word983 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X355 GND A5 word714 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X356 a_710_n8010# A7 a_446_n8010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X357 a_1898_n48906# a_1848_n66# a_1766_n48906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X358 word53 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X359 a_446_n97186# A8 a_50_n97186# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X360 a_2030_n7442# A2 a_1766_n7442# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X361 a_842_n15110# a_792_n66# a_710_n15110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X362 word491 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X363 word222 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X364 a_974_n44646# A6 a_710_n44646# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X365 GND A6 word401 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X366 GND A3 word1014 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X367 word95 a_2376_n66# a_2162_n13690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X368 word938 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X369 word803 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X370 word744 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X371 a_710_n7584# A7 a_446_n7584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X372 a_842_n84406# a_792_n66# a_710_n84406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X373 GND A8 word585 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X374 word919 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X375 a_50_n109540# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X376 word583 a_2376_n66# a_2162_n82986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X377 GND A2 word906 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X378 a_842_n14684# a_792_n66# a_710_n14684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X379 a_50_n131976# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X380 a_50_n140354# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X381 word434 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X382 GND A4 word396 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X383 word427 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X384 a_1106_n51178# a_1056_n66# a_842_n51178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X385 word967 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X386 a_578_n34848# a_528_n66# a_446_n34848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X387 a_1106_n42800# a_1056_n66# a_974_n42800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X388 a_842_n123314# a_792_n66# a_710_n123314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X389 a_50_n117492# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X390 a_1898_n16956# a_1848_n66# a_1766_n16956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X391 word273 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X392 a_1106_n98038# a_1056_n66# a_974_n98038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X393 a_182_n64952# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X394 a_314_n126722# a_264_n66# a_50_n126722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X395 a_1106_n89660# a_1056_n66# a_842_n89660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X396 a_974_n21074# A6 a_578_n21074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X397 word1010 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X398 word266 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X399 a_2030_n484# A2 a_1766_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X400 a_1502_n6732# A4 a_1106_n6732# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X401 GND A6 word176 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X402 a_50_n73472# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X403 a_842_n52456# a_792_n66# a_710_n52456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X404 word327 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X405 a_974_n59556# A6 a_578_n59556# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X406 GND A0 word610 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X407 a_182_n33428# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X408 GND A0 word178 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X409 a_182_n6874# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X410 a_314_n71342# a_264_n66# a_182_n71342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X411 a_1502_n15536# A4 a_1106_n15536# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X412 a_1370_n98890# a_1320_n66# a_1106_n98890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X413 GND A8 word690 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X414 a_314_n62964# a_264_n66# a_182_n62964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X415 word167 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X416 GND A4 word171 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X417 a_842_n29594# a_792_n66# a_578_n29594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X418 a_578_n72620# a_528_n66# a_314_n72620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X419 word598 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X420 word539 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X421 GND A0 word666 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X422 word742 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X423 word834 A0 a_2162_n118628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X424 a_2030_n4886# A2 a_1766_n4886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X425 a_578_n58136# a_528_n66# a_314_n58136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X426 a_842_n138224# a_792_n66# a_578_n138224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X427 a_1370_n7442# a_1320_n66# a_1106_n7442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X428 GND A3 word341 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X429 GND A4 word13 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X430 a_842_n90228# a_792_n66# a_710_n90228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X431 a_974_n97328# A6 a_578_n97328# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X432 word102 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X433 a_1634_n17524# a_1584_n66# a_1370_n17524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X434 GND A0 word444 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X435 GND A2 word947 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X436 word7 a_2376_n66# a_2162_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X437 word656 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X438 word597 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X439 word310 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X440 a_50_n88382# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X441 a_842_n67366# a_792_n66# a_578_n67366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X442 word163 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X443 word949 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X444 a_842_n120758# a_792_n66# a_710_n120758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X445 a_182_n48338# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X446 a_1898_n5596# a_1848_n66# a_1766_n5596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X447 a_1898_n22778# a_1848_n66# a_1634_n22778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X448 word314 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X449 word373 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X450 a_182_n39960# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X451 a_182_n70774# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X452 word331 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X453 word336 A0 a_2294_n47912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X454 a_314_n132544# a_264_n66# a_50_n132544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X455 a_1898_n78016# a_1848_n66# a_1766_n78016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X456 GND A6 word649 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X457 word651 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X458 word366 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X459 a_1106_n135952# a_1056_n66# a_974_n135952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X460 word143 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X461 word307 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X462 a_578_n26186# a_528_n66# a_446_n26186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X463 a_842_n106274# a_792_n66# a_578_n106274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X464 a_1766_n136804# A3 a_1502_n136804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X465 GND A3 word116 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X466 GND A8 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X467 a_1634_n46918# a_1584_n66# a_1502_n46918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X468 a_974_n57000# A6 a_578_n57000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X469 a_314_n109682# a_264_n66# a_50_n109682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X470 word890 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X471 a_314_n46350# a_264_n66# a_182_n46350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X472 a_578_n95482# a_528_n66# a_446_n95482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X473 GND A4 word644 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X474 GND A2 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X475 word429 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X476 word930 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X477 word207 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X478 GND A0 word490 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X479 a_1502_n59840# A4 a_1106_n59840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X480 word415 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X481 word783 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X482 GND A4 word483 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X483 word702 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X484 a_182_n16388# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X485 word860 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X486 word106 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X487 word209 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X488 a_842_n144046# a_792_n66# a_578_n144046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X489 a_578_n55580# a_528_n66# a_314_n55580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X490 word478 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X491 word426 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X492 a_2294_n44504# A1 a_2030_n44504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X493 word108 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X494 word575 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X495 a_1766_n104854# A3 a_1502_n104854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X496 word471 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X497 GND A6 word695 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X498 a_710_n41522# A7 a_314_n41522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X499 a_1634_n14968# a_1584_n66# a_1502_n14968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X500 word916 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X501 word857 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X502 word638 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X503 word722 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X504 a_1898_n113516# a_1848_n66# a_1634_n113516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X505 word414 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X506 word145 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X507 word596 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X508 word990 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X509 a_1634_n92642# a_1584_n66# a_1502_n92642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X510 a_182_n54160# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X511 word436 A0 a_2294_n62112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X512 a_1502_n27890# A4 a_1238_n27890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X513 word475 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X514 a_1634_n142342# a_1584_n66# a_1502_n142342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X515 a_1106_n141774# a_1056_n66# a_842_n141774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X516 a_1634_n133964# a_1584_n66# a_1502_n133964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X517 word980 A0 a_2294_n139360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X518 word306 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X519 a_1238_n13548# A5 a_842_n13548# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X520 word374 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X521 GND A6 word927 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X522 GND A9 word91 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X523 word965 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X524 a_974_n130840# A6 a_578_n130840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X525 a_1634_n61118# a_1584_n66# a_1502_n61118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X526 word455 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X527 GND A5 word586 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X528 a_2030_n121752# A2 a_1634_n121752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X529 GND A3 word487 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X530 a_1238_n82844# A5 a_842_n82844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X531 a_1238_n91222# A5 a_974_n91222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X532 a_1898_n142910# a_1848_n66# a_1634_n142910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X533 a_2162_n52314# a_2112_n66# a_1898_n52314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X534 a_2294_n59414# A1 a_2030_n59414# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X535 a_1766_n128142# A3 a_1502_n128142# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X536 a_974_n116356# A6 a_710_n116356# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X537 a_1634_n38256# a_1584_n66# a_1502_n38256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X538 word371 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X539 a_1502_n74040# A4 a_1238_n74040# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X540 word1021 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X541 a_1634_n60692# a_1584_n66# a_1502_n60692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X542 word511 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X543 word886 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X544 word59 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X545 word579 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X546 a_1898_n128426# a_1848_n66# a_1766_n128426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X547 a_2162_n114652# a_2112_n66# a_1898_n114652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X548 word152 A0 a_2294_n21784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X549 a_842_n88098# a_792_n66# a_710_n88098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X550 word147 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X551 a_2162_n29452# a_2112_n66# a_1898_n29452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X552 word250 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X553 a_1634_n110392# a_1584_n66# a_1502_n110392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X554 a_446_n33712# A8 a_182_n33712# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X555 word572 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X556 GND A7 word829 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X557 a_842_n141490# a_792_n66# a_578_n141490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X558 a_182_n69070# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X559 GND A3 word423 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X560 word482 A0 a_2162_n68644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X561 GND A9 word298 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X562 a_2030_n128710# A2 a_1634_n128710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X563 a_2294_n50326# A1 a_2030_n50326# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X564 word891 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X565 word418 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X566 a_314_n144898# a_264_n66# a_50_n144898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X567 a_710_n16530# A7 a_446_n16530# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X568 word90 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X569 GND A5 word203 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X570 word289 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X571 word740 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X572 a_2294_n118912# A1 a_1898_n118912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X573 GND A3 word694 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X574 a_1238_n28458# A5 a_842_n28458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X575 a_2162_n81708# a_2112_n66# a_1898_n81708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X576 a_2294_n88808# A1 a_2030_n88808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X577 word479 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X578 GND A9 word196 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X579 a_2030_n76312# A2 a_1634_n76312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X580 GND A9 word137 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X581 a_2030_n136662# A2 a_1766_n136662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X582 a_1898_n110960# a_1848_n66# a_1634_n110960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X583 a_2162_n20364# a_2112_n66# a_1898_n20364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X584 a_2294_n27464# A1 a_2030_n27464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X585 a_1634_n67650# a_1584_n66# a_1370_n67650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X586 a_710_n85826# A7 a_446_n85826# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X587 word637 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X588 a_2162_n11986# a_2112_n66# a_2030_n11986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X589 word260 A0 a_2294_n37120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X590 a_1502_n42090# A4 a_1106_n42090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X591 word946 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X592 a_1106_n125160# a_1056_n66# a_842_n125160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X593 a_1634_n117350# a_1584_n66# a_1370_n117350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X594 word354 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X595 word189 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X596 word476 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X597 GND A6 word810 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X598 GND A5 word80 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X599 GND A9 word505 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X600 a_2162_n129562# a_2112_n66# a_1898_n129562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X601 word316 A0 a_2294_n45072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X602 a_2030_n105138# A2 a_1766_n105138# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X603 GND A9 word73 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X604 GND A5 word410 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X605 word677 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X606 a_1238_n66230# A5 a_842_n66230# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X607 word618 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X608 word724 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X609 GND A3 word528 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X610 GND A9 word403 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X611 GND A3 word469 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X612 GND A6 word807 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X613 word195 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X614 word254 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X615 word731 a_2376_n66# a_2162_n104002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X616 a_1766_n125586# A3 a_1370_n125586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X617 a_974_n113800# A6 a_710_n113800# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X618 word335 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X619 a_1634_n35700# a_1584_n66# a_1370_n35700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X620 a_710_n53876# A7 a_314_n53876# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X621 GND A5 word407 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X622 GND A5 word466 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X623 word868 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X624 a_1238_n74182# A5 a_974_n74182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X625 GND A8 word243 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X626 a_2162_n96618# a_2112_n66# a_1898_n96618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X627 a_1238_n139502# A5 a_842_n139502# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X628 a_2162_n120474# a_2112_n66# a_1898_n120474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X629 word721 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X630 a_1898_n125870# a_1848_n66# a_1766_n125870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X631 a_2162_n35274# a_2112_n66# a_1898_n35274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X632 GND A7 word96 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X633 a_710_n39392# A7 a_314_n39392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X634 a_1766_n21642# A3 a_1370_n21642# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X635 GND A1 word236 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X636 GND A7 word870 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X637 GND A9 word11 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X638 GND A0 word836 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X639 word459 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X640 a_1766_n68502# A3 a_1502_n68502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X641 a_2294_n133112# A1 a_2030_n133112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X642 a_2294_n124734# A1 a_1898_n124734# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X643 a_446_n16672# A8 a_182_n16672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X644 word89 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X645 GND A7 word768 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X646 GND A1 word993 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X647 a_1106_n7016# a_1056_n66# a_974_n7016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X648 a_2294_n94630# A1 a_2030_n94630# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X649 word862 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X650 a_1238_n130414# A5 a_974_n130414# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X651 a_2030_n82134# A2 a_1766_n82134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X652 GND A9 word178 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X653 a_2030_n142484# A2 a_1634_n142484# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X654 word771 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X655 a_2294_n33286# A1 a_2030_n33286# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X656 a_578_n135952# a_528_n66# a_314_n135952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X657 word26 A0 a_2162_n3892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X658 word169 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X659 word636 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X660 a_1370_n11844# a_1320_n66# a_1238_n11844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X661 word987 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X662 GND A8 word77 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X663 GND A7 word362 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X664 word928 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X665 GND A1 word832 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X666 GND A1 word773 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X667 a_2162_n64668# a_2112_n66# a_1898_n64668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X668 a_446_n104144# A8 a_50_n104144# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X669 a_1898_n102298# a_1848_n66# a_1634_n102298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X670 GND A9 word60 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X671 a_1370_n58704# a_1320_n66# a_1238_n58704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X672 a_710_n77164# A7 a_446_n77164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X673 a_2030_n59272# A2 a_1766_n59272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X674 GND A6 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X675 word657 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X676 word973 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X677 a_1370_n116214# a_1320_n66# a_1106_n116214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X678 a_578_n104428# a_528_n66# a_446_n104428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X679 a_1370_n107836# a_1320_n66# a_1106_n107836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X680 GND A1 word341 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X681 word707 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X682 a_1766_n36552# A3 a_1502_n36552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X683 word628 A0 a_2294_n89376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X684 GND A9 word444 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X685 a_1106_n17524# a_1056_n66# a_842_n17524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X686 GND A4 word998 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X687 GND A9 word385 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X688 a_2294_n62680# A1 a_2030_n62680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X689 GND A1 word709 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X690 word253 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X691 a_2030_n50184# A2 a_1766_n50184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X692 word713 a_2376_n66# a_2294_n101446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X693 a_1238_n49190# A5 a_842_n49190# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X694 word557 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X695 word715 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X696 word850 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X697 word967 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X698 a_1238_n136946# A5 a_842_n136946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X699 a_2030_n97044# A2 a_1634_n97044# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X700 GND A4 word896 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X701 a_710_n121042# A7 a_314_n121042# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X702 GND A6 word55 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X703 a_710_n112664# A7 a_314_n112664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X704 a_1370_n35132# a_1320_n66# a_1106_n35132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X705 GND A8 word21 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X706 word948 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X707 GND A0 word936 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X708 a_1370_n26754# a_1320_n66# a_1106_n26754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X709 GND A8 word182 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X710 word564 A0 a_2294_n80288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X711 GND A8 word123 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X712 a_2162_n79578# a_2112_n66# a_1898_n79578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X713 a_2294_n108120# A1 a_2030_n108120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X714 a_446_n83838# A8 a_50_n83838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X715 a_446_n92216# A8 a_50_n92216# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X716 a_446_n22494# A8 a_182_n22494# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X717 GND A1 word116 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X718 GND A6 word52 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X719 GND A7 word809 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X720 GND A2 word184 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X721 GND A8 word611 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X722 GND A9 word219 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X723 word460 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X724 a_2294_n116072# A1 a_2030_n116072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X725 a_578_n141774# a_528_n66# a_314_n141774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X726 a_710_n2614# A7 a_446_n2614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X727 a_2294_n107694# A1 a_1898_n107694# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X728 GND A2 word672 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X729 GND A9 word490 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X730 a_2294_n77590# A1 a_2030_n77590# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X731 GND A1 word873 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X732 GND A3 word818 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X733 a_1238_n113374# A5 a_974_n113374# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X734 a_2162_n70490# a_2112_n66# a_1898_n70490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X735 a_446_n101588# A8 a_50_n101588# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X736 GND A3 word759 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X737 a_2030_n65094# A2 a_1634_n65094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X738 word759 a_2376_n66# a_2162_n107978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X739 word1014 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X740 word879 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X741 a_1370_n122036# a_1320_n66# a_1238_n122036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X742 word723 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X743 a_1370_n113658# a_1320_n66# a_1238_n113658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X744 a_50_n112522# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X745 GND A5 word784 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X746 word7 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X747 GND A0 word982 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X748 a_1106_n23346# a_1056_n66# a_974_n23346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X749 GND A6 word141 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X750 a_1766_n89234# A3 a_1370_n89234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X751 word1019 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X752 a_1106_n14968# a_1056_n66# a_842_n14968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X753 a_446_n98748# A8 a_50_n98748# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X754 word876 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X755 word235 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X756 word165 a_2376_n66# a_2294_n23630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X757 GND A6 word412 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X758 word949 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X759 word1008 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X760 GND A2 word506 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X761 GND A4 word937 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X762 GND A4 word878 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X763 a_182_n1904# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X764 a_1370_n93920# a_1320_n66# a_1238_n93920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X765 a_2030_n94488# A2 a_1634_n94488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X766 GND A8 word655 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X767 GND A0 word760 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X768 word989 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X769 a_842_n33002# a_792_n66# a_578_n33002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X770 GND A8 word725 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X771 GND A0 word918 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X772 a_2162_n9146# a_2112_n66# a_1898_n9146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X773 GND A8 word164 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X774 GND A1 word648 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X775 word653 a_2376_n66# a_2294_n92926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X776 a_1238_n128284# A5 a_974_n128284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X777 a_50_n141916# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X778 word221 a_2376_n66# a_2294_n31582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X779 a_1766_n80146# A3 a_1370_n80146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X780 GND A1 word589 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X781 GND A1 word157 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X782 a_1106_n61118# a_1056_n66# a_974_n61118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X783 word621 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X784 word887 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X785 word828 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X786 a_1370_n18092# a_1320_n66# a_1106_n18092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X787 GND A2 word225 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X788 a_1106_n52740# a_1056_n66# a_842_n52740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X789 word551 a_2376_n66# a_2162_n78442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X790 GND A8 word652 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X791 GND A0 word816 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X792 a_446_n4034# A8 a_182_n4034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X793 a_50_n127432# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X794 GND A7 word347 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X795 a_446_n75176# A8 a_50_n75176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X796 word343 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X797 a_1766_n57284# A3 a_1370_n57284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X798 GND A2 word555 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X799 word336 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X800 a_1502_n137230# A4 a_1238_n137230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X801 a_974_n22636# A6 a_578_n22636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X802 GND A6 word187 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X803 a_1106_n60692# a_1056_n66# a_974_n60692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X804 word783 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X805 word859 a_2376_n66# a_2162_n122178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X806 GND A3 word800 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X807 a_50_n83412# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X808 a_1370_n61970# a_1320_n66# a_1106_n61970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X809 a_2294_n6022# A1 a_2030_n6022# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X810 a_974_n91932# A6 a_578_n91932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X811 word5 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X812 GND A0 word248 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X813 GND A7 word283 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X814 GND A2 word552 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X815 a_974_n2188# A6 a_710_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X816 GND A1 word364 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X817 GND A7 word613 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X818 GND A7 word554 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X819 word812 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X820 a_3292_164# A1 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X821 a_578_n21216# a_528_n66# a_446_n21216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X822 a_1766_n86678# A3 a_1502_n86678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X823 a_842_n101304# a_792_n66# a_578_n101304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X824 GND A5 word20 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X825 word118 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X826 word177 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X827 a_182_n42942# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X828 GND A3 word81 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X829 a_974_n60408# A6 a_578_n60408# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X830 GND A2 word330 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X831 a_1502_n105280# A4 a_1106_n105280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X832 word990 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X833 word62 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X834 a_974_n37546# A6 a_710_n37546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X835 word231 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X836 a_842_n30446# a_792_n66# a_578_n30446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X837 word172 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X838 GND A2 word1017 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X839 word888 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X840 GND A3 word964 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X841 word667 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X842 word753 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X843 a_182_n11418# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X844 a_50_n98322# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X845 GND A4 word448 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X846 a_1370_n85258# a_1320_n66# a_1238_n85258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X847 a_314_n40954# a_264_n66# a_182_n40954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X848 a_50_n89944# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X849 a_842_n68928# a_792_n66# a_578_n68928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X850 a_1370_n76880# a_1320_n66# a_1238_n76880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X851 GND A8 word535 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X852 word174 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X853 word734 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X854 a_1370_n134390# a_1320_n66# a_1106_n134390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X855 a_50_n133254# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X856 a_1898_n32718# a_1848_n66# a_1766_n32718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X857 word443 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X858 word533 a_2376_n66# a_2294_n75886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X859 a_446_n1478# A8 a_182_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X860 a_50_n124876# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X861 GND A1 word469 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X862 GND A1 word528 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X863 word436 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X864 GND A6 word660 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X865 word377 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X866 a_182_n10992# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X867 a_578_n36126# a_528_n66# a_446_n36126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X868 a_1238_n9714# A5 a_842_n9714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X869 a_1106_n35700# a_1056_n66# a_842_n35700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X870 a_1106_n44078# a_1056_n66# a_974_n44078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X871 a_578_n27748# a_528_n66# a_446_n27748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X872 a_1898_n18234# a_1848_n66# a_1634_n18234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X873 a_842_n107836# a_792_n66# a_578_n107836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X874 word29 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X875 a_182_n57852# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X876 a_50_n80856# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X877 a_974_n75318# A6 a_710_n75318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X878 a_314_n119622# a_264_n66# a_50_n119622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X879 GND A5 word769 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X880 a_1634_n2046# a_1584_n66# a_1502_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X881 GND A6 word558 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X882 GND A0 word230 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X883 GND A2 word851 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X884 GND A2 word792 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X885 a_1502_n22920# A4 a_1106_n22920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X886 word277 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X887 GND A0 word560 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X888 word26 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X889 GND A7 word595 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X890 word853 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X891 a_1766_n7868# A3 a_1370_n7868# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X892 GND A0 word128 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X893 a_974_n74892# A6 a_710_n74892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X894 GND A4 word612 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X895 a_182_n8152# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X896 a_182_n26328# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X897 word159 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X898 word218 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X899 GND A4 word553 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X900 word1016 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X901 a_182_n17950# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X902 a_314_n55864# a_264_n66# a_182_n55864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X903 a_314_n64242# a_264_n66# a_182_n64242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X904 a_1106_n113942# a_1056_n66# a_974_n113942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X905 a_578_n65520# a_528_n66# a_314_n65520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X906 a_1898_n47628# a_1848_n66# a_1634_n47628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X907 a_314_n110534# a_264_n66# a_50_n110534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X908 word697 a_2376_n66# a_2294_n99174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X909 word496 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X910 word839 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X911 GND A6 word435 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X912 GND A0 word616 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X913 a_50_n139786# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X914 a_2030_n6164# A2 a_1634_n6164# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X915 GND A3 word34 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X916 word44 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X917 a_1502_n77732# A4 a_1106_n77732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X918 word482 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X919 word942 A0 a_2162_n133964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X920 a_974_n43368# A6 a_710_n43368# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X921 a_1634_n24908# a_1584_n66# a_1502_n24908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X922 word213 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X923 word986 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X924 word927 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X925 word543 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X926 a_50_n95766# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X927 GND A4 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X928 word484 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X929 a_842_n83128# a_792_n66# a_710_n83128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X930 GND A0 word394 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X931 word215 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X932 word633 a_2376_n66# a_2294_n90086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X933 word775 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X934 a_1634_n8578# a_1584_n66# a_1370_n8578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X935 a_2294_n9998# A1 a_1898_n9998# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X936 a_1502_n46208# A4 a_1238_n46208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X937 word720 A0 a_2294_n102440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X938 GND A2 word897 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X939 a_50_n130698# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X940 a_1502_n37830# A4 a_1238_n37830# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X941 word547 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X942 word606 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X943 word766 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X944 word260 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X945 GND A4 word328 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X946 GND A4 word387 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X947 word705 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X948 word958 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X949 a_842_n122036# a_792_n66# a_710_n122036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X950 a_578_n33570# a_528_n66# a_446_n33570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X951 a_1898_n15678# a_1848_n66# a_1634_n15678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X952 a_182_n72052# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X953 GND A3 word227 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X954 a_182_n63674# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X955 a_1502_n45782# A4 a_1238_n45782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X956 a_974_n81140# A6 a_710_n81140# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X957 a_314_n125444# a_264_n66# a_50_n125444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X958 word776 A0 a_2294_n110392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X959 GND A6 word540 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X960 word316 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X961 word257 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X962 word93 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X963 a_578_n19086# a_528_n66# a_446_n19086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X964 a_1502_n5454# A4 a_1106_n5454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X965 a_1898_n84974# a_1848_n66# a_1766_n84974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X966 a_1766_n129704# A3 a_1370_n129704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X967 a_842_n51178# a_792_n66# a_710_n51178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X968 a_974_n58278# A6 a_578_n58278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X969 word318 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X970 a_974_n117918# A6 a_710_n117918# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X971 word581 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X972 a_182_n5596# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X973 a_182_n32150# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X974 a_314_n39250# a_264_n66# a_182_n39250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X975 a_314_n70064# a_264_n66# a_182_n70064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X976 a_1502_n14258# A4 a_1106_n14258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X977 word222 A0 a_2162_n31724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X978 a_314_n61686# a_264_n66# a_182_n61686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X979 a_842_n89660# a_792_n66# a_710_n89660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X980 a_1634_n120332# a_1584_n66# a_1502_n120332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X981 word158 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X982 a_1898_n53450# a_1848_n66# a_1766_n53450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X983 word530 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X984 word733 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X985 GND A3 word434 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X986 a_1502_n83554# A4 a_1238_n83554# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X987 GND A0 word48 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X988 a_1766_n120616# A3 a_1370_n120616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X989 word646 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X990 word810 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X991 word481 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X992 a_974_n96050# A6 a_578_n96050# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X993 GND A3 word273 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X994 word525 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X995 word139 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X996 a_1502_n52030# A4 a_1106_n52030# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X997 word216 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X998 a_1898_n99884# a_1848_n66# a_1634_n99884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X999 word866 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1000 GND A2 word938 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1001 word588 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1002 word807 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1003 word647 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1004 word731 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1005 a_1898_n106416# a_1848_n66# a_1634_n106416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1006 a_1238_n37972# A5 a_974_n37972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1007 a_842_n66088# a_792_n66# a_578_n66088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1008 word154 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1009 word999 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1010 a_1634_n85542# a_1584_n66# a_1370_n85542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1011 word940 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1012 a_446_n11702# A8 a_182_n11702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1013 a_1898_n21500# a_1848_n66# a_1766_n21500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1014 word386 A0 a_2162_n55012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1015 a_182_n47060# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1016 a_1502_n29168# A4 a_1238_n29168# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1017 GND A9 word143 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1018 a_1106_n143052# a_1056_n66# a_842_n143052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1019 a_314_n131266# a_264_n66# a_50_n131266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1020 GND A6 word640 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1021 a_1106_n134674# a_1056_n66# a_974_n134674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1022 a_1634_n126864# a_1584_n66# a_1370_n126864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1023 word263 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1024 a_314_n122888# a_264_n66# a_50_n122888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1025 word642 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1026 word75 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1027 GND A3 word598 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1028 GND A6 word936 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1029 word838 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1030 a_1898_n90796# a_1848_n66# a_1634_n90796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1031 word324 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1032 a_974_n132118# A6 a_578_n132118# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1033 word359 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1034 a_1634_n54018# a_1584_n66# a_1370_n54018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1035 word405 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1036 word300 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1037 a_2030_n45924# A2 a_1766_n45924# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1038 GND A5 word536 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1039 GND A5 word477 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1040 a_1238_n84122# A5 a_842_n84122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1041 a_1502_n20080# A4 a_1238_n20080# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1042 a_1238_n75744# A5 a_974_n75744# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1043 word630 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1044 a_974_n109256# A6 a_710_n109256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1045 a_2162_n36836# a_2112_n66# a_2030_n36836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1046 a_710_n49332# A7 a_314_n49332# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1047 word321 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1048 word971 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1049 a_974_n131692# A6 a_578_n131692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1050 a_1634_n53592# a_1584_n66# a_1370_n53592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1051 word461 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1052 GND A0 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1053 word470 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1054 GND A0 word30 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1055 word102 A0 a_2162_n14684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1056 a_446_n26612# A8 a_182_n26612# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1057 word200 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1058 GND A3 word373 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1059 GND A9 word248 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1060 a_314_n137798# a_264_n66# a_50_n137798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1061 word841 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1062 a_2294_n34848# A1 a_1898_n34848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1063 word99 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1064 word688 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1065 a_1634_n13690# a_1584_n66# a_1370_n13690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1066 a_710_n40244# A7 a_314_n40244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1067 a_1634_n22068# a_1584_n66# a_1370_n22068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1068 word239 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1069 word526 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1070 a_2030_n13974# A2 a_1766_n13974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1071 word998 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1072 word713 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1073 a_446_n105706# A8 a_50_n105706# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1074 a_1898_n112238# a_1848_n66# a_1766_n112238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1075 a_710_n78726# A7 a_446_n78726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1076 a_710_n87104# A7 a_446_n87104# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1077 word587 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1078 GND A1 word81 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1079 a_710_n17382# A7 a_446_n17382# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1080 GND A6 word17 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1081 GND A7 word774 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1082 word984 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1083 a_2162_n145324# a_2112_n66# a_1898_n145324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1084 a_2162_n136946# a_2112_n66# a_2030_n136946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1085 word368 A0 a_2294_n52456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1086 word896 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1087 a_1106_n118060# a_1056_n66# a_974_n118060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1088 word777 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1089 a_2294_n111102# A1 a_1898_n111102# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1090 word698 A0 a_2162_n99316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1091 a_1238_n12270# A5 a_842_n12270# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1092 word238 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1093 word297 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1094 GND A3 word580 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1095 GND A6 word918 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1096 GND A9 word455 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1097 word365 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1098 a_1766_n141348# A3 a_1502_n141348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1099 a_1766_n132970# A3 a_1502_n132970# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1100 GND A2 word146 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1101 a_2030_n51746# A2 a_1634_n51746# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1102 a_1238_n59130# A5 a_974_n59130# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1103 GND A5 word577 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1104 word627 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1105 GND A5 word518 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1106 GND A3 word419 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1107 GND A6 word816 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1108 a_2294_n49758# A1 a_1898_n49758# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1109 a_2162_n51036# a_2112_n66# a_1898_n51036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1110 word204 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1111 a_2294_n58136# A1 a_2030_n58136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1112 GND A9 word511 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1113 a_1766_n118486# A3 a_1502_n118486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1114 a_710_n122604# A7 a_314_n122604# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1115 a_974_n115078# A6 a_710_n115078# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1116 a_2162_n42658# a_2112_n66# a_2030_n42658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1117 a_1634_n28600# a_1584_n66# a_1502_n28600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1118 a_2030_n28884# A2 a_1634_n28884# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1119 a_710_n46776# A7 a_314_n46776# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1120 GND A8 word32 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1121 word634 A0 a_2162_n90228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1122 word50 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1123 GND A8 word193 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1124 word759 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1125 a_1238_n67082# A5 a_842_n67082# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1126 word570 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1127 a_2162_n104996# a_2112_n66# a_2030_n104996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1128 a_1898_n127148# a_1848_n66# a_1634_n127148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1129 a_842_n9430# a_792_n66# a_710_n9430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1130 a_446_n32434# A8 a_182_n32434# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1131 a_1766_n14542# A3 a_1502_n14542# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1132 a_2162_n19796# a_2112_n66# a_2030_n19796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1133 word563 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1134 GND A7 word879 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1135 word504 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1136 GND A7 word820 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1137 word414 A0 a_2162_n58988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1138 GND A8 word681 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1139 GND A9 word289 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1140 GND A9 word230 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1141 GND A8 word751 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1142 a_2294_n40670# A1 a_1898_n40670# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1143 word350 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1144 GND A5 word135 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1145 GND A7 word51 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1146 GND A7 word876 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1147 word812 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1148 GND A9 word128 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1149 GND A1 word884 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1150 GND A2 word251 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1151 a_710_n84548# A7 a_446_n84548# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1152 a_2030_n135384# A2 a_1634_n135384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1153 word829 a_2376_n66# a_2294_n117918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1154 a_578_n128852# a_528_n66# a_314_n128852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1155 GND A4 word741 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1156 a_1370_n13122# a_1320_n66# a_1238_n13122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1157 word119 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1158 word586 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1159 word793 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1160 GND A0 word722 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1161 word937 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1162 GND A7 word312 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1163 a_974_n6306# A6 a_710_n6306# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1164 a_1766_n43936# A3 a_1370_n43936# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1165 word607 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1166 word680 A0 a_2294_n96760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1167 word675 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1168 a_2162_n128284# a_2112_n66# a_1898_n128284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1169 a_1106_n24908# a_1056_n66# a_974_n24908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1170 a_1370_n109114# a_1320_n66# a_1106_n109114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1171 word609 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1172 GND A9 word394 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1173 GND A9 word66 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1174 GND A9 word335 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1175 word203 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1176 a_710_n52598# A7 a_314_n52598# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1177 GND A5 word457 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1178 word361 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1179 GND A8 word234 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1180 a_2162_n95340# a_2112_n66# a_1898_n95340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1181 word859 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1182 a_1238_n138224# A5 a_842_n138224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1183 a_1370_n100026# a_1320_n66# a_1106_n100026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1184 a_1238_n129846# A5 a_974_n129846# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1185 GND A7 word87 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1186 word291 a_2376_n66# a_2162_n41522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1187 a_1766_n11986# A3 a_1370_n11986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1188 word632 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1189 GND A0 word886 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1190 a_446_n910# A8 a_182_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1191 word514 A0 a_2162_n73188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1192 a_1502_n100310# A4 a_1238_n100310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1193 word983 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1194 word20 A0 a_2294_n3040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1195 a_446_n85116# A8 a_50_n85116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1196 word450 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1197 word923 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1198 a_446_n76738# A8 a_50_n76738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1199 a_2294_n123456# A1 a_1898_n123456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1200 a_446_n15394# A8 a_182_n15394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1201 GND A3 word929 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1202 a_2162_n1620# a_2112_n66# a_2030_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1203 GND A7 word33 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1204 a_1106_n70632# a_1056_n66# a_842_n70632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1205 word794 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1206 word853 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1207 GND A8 word561 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1208 GND A9 word169 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1209 word929 a_2376_n66# a_2294_n132118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1210 GND A1 word925 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1211 GND A3 word870 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1212 a_1238_n120758# A5 a_842_n120758# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1213 a_710_n90370# A7 a_446_n90370# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1214 GND A4 word782 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1215 a_578_n143052# a_528_n66# a_314_n143052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1216 a_578_n134674# a_528_n66# a_314_n134674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1217 word410 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1218 a_1370_n71910# a_1320_n66# a_1106_n71910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1219 GND A5 word664 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1220 word51 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1221 word568 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1222 GND A7 word353 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1223 word919 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1224 GND A1 word493 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1225 GND A7 word294 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1226 GND A3 word768 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1227 GND A1 word764 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1228 a_974_n3750# A6 a_710_n3750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1229 a_1370_n57426# a_1320_n66# a_1238_n57426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1230 word964 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1231 GND A7 word624 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1232 word732 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1233 a_578_n103150# a_528_n66# a_446_n103150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1234 a_1766_n96618# A3 a_1502_n96618# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1235 a_50_n105422# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1236 word987 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1237 a_1766_n35274# A3 a_1370_n35274# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1238 GND A1 word273 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1239 GND A1 word332 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1240 GND A5 word734 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1241 a_1502_n115220# A4 a_1106_n115220# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1242 a_1106_n16246# a_1056_n66# a_842_n16246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1243 GND A3 word704 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1244 word969 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1245 a_2294_n138366# A1 a_1898_n138366# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1246 word826 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1247 GND A1 word57 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1248 word185 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1249 word958 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1250 word115 a_2376_n66# a_2162_n16530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1251 word899 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1252 a_710_n111386# A7 a_314_n111386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1253 word975 a_2376_n66# a_2162_n138650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1254 a_1502_n123172# A4 a_1106_n123172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1255 a_1502_n114794# A4 a_1106_n114794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1256 GND A8 word605 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1257 a_182_n200# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1258 a_1370_n144330# a_1320_n66# a_1106_n144330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1259 a_842_n17524# a_792_n66# a_710_n17524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1260 a_1370_n25476# a_1320_n66# a_1106_n25476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1261 word603 a_2376_n66# a_2162_n85826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1262 GND A0 word868 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1263 a_50_n134816# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1264 a_1766_n73046# A3 a_1502_n73046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1265 GND A8 word114 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1266 a_2162_n78300# a_2112_n66# a_1898_n78300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1267 word171 a_2376_n66# a_2162_n24482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1268 a_446_n82560# A8 a_50_n82560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1269 a_1766_n64668# A3 a_1502_n64668# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1270 a_182_n20932# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1271 a_1106_n54018# a_1056_n66# a_842_n54018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1272 a_1370_n94772# a_1320_n66# a_1238_n94772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1273 GND A8 word661 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1274 GND A6 word298 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1275 GND A8 word602 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1276 a_578_n140496# a_528_n66# a_314_n140496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1277 a_710_n1336# A7 a_446_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1278 GND A5 word839 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1279 a_1634_n3608# a_1584_n66# a_1370_n3608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1280 GND A6 word137 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1281 GND A9 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1282 a_1238_n112096# A5 a_974_n112096# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1283 a_1106_n53592# a_1056_n66# a_842_n53592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1284 word512 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1285 word809 a_2376_n66# a_2294_n115078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1286 a_50_n76312# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1287 GND A4 word293 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1288 a_1370_n63248# a_1320_n66# a_1106_n63248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1289 a_842_n46918# a_792_n66# a_710_n46918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1290 word507 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1291 GND A0 word198 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1292 word437 a_2376_n66# a_2294_n62254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1293 a_1502_n138082# A4 a_1238_n138082# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1294 a_1370_n112380# a_1320_n66# a_1238_n112380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1295 a_182_n9714# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1296 a_50_n111244# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1297 a_710_n126296# A7 a_314_n126296# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1298 a_314_n65804# a_264_n66# a_182_n65804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1299 a_50_n102866# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1300 a_1766_n41096# A3 a_1502_n41096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1301 GND A0 word356 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1302 GND A1 word373 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1303 GND A4 word132 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1304 word281 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1305 GND A5 word775 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1306 GND A0 word914 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1307 a_446_n97470# A8 a_50_n97470# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1308 GND A0 word686 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1309 word127 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1310 word1012 A0 a_2294_n143904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1311 a_182_n35842# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1312 a_974_n44930# A6 a_710_n44930# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1313 GND A6 word403 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1314 word999 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1315 word940 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1316 word906 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1317 GND A4 word869 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1318 word805 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1319 a_710_n7868# A7 a_446_n7868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1320 word27 a_2376_n66# a_2162_n4034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1321 a_1370_n31298# a_1320_n66# a_1238_n31298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1322 GND A0 word850 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1323 a_842_n14968# a_792_n66# a_710_n14968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1324 a_50_n140638# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1325 word838 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1326 word836 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1327 GND A4 word398 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1328 GND A1 word580 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1329 word617 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1330 a_314_n42232# a_264_n66# a_182_n42232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1331 a_974_n99742# A6 a_578_n99742# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1332 word819 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1333 word483 a_2376_n66# a_2162_n68786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1334 GND A7 word338 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1335 a_1370_n127290# a_1320_n66# a_1106_n127290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1336 a_50_n117776# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1337 a_50_n126154# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1338 a_1502_n55722# A4 a_1238_n55722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1339 word846 A0 a_2162_n120332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1340 word386 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1341 word327 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1342 a_974_n21358# A6 a_578_n21358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1343 a_578_n29026# a_528_n66# a_446_n29026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1344 GND A6 word178 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1345 a_842_n109114# a_792_n66# a_578_n109114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1346 a_50_n82134# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1347 a_50_n73756# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1348 a_842_n52740# a_792_n66# a_710_n52740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1349 a_974_n59840# A6 a_578_n59840# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1350 a_578_n98322# a_528_n66# a_446_n98322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1351 a_1106_n97896# a_1056_n66# a_974_n97896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1352 GND A0 word180 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1353 GND A6 word666 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1354 a_314_n71626# a_264_n66# a_182_n71626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1355 a_1502_n15820# A4 a_1106_n15820# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1356 GND A4 word173 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1357 GND A4 word232 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1358 GND A0 word1014 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1359 GND A7 word545 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1360 a_842_n29878# a_792_n66# a_578_n29878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1361 GND A1 word685 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1362 a_182_n19228# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1363 a_182_n50042# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1364 a_314_n57142# a_264_n66# a_182_n57142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1365 a_182_n41664# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1366 a_314_n48764# a_264_n66# a_182_n48764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1367 a_1502_n23772# A4 a_1106_n23772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1368 GND A6 word444 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1369 a_1106_n106842# a_1056_n66# a_842_n106842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1370 a_1370_n7726# a_1320_n66# a_1106_n7726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1371 a_578_n58420# a_528_n66# a_314_n58420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1372 GND A6 word385 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1373 word446 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1374 word1006 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1375 a_842_n138508# a_792_n66# a_578_n138508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1376 a_446_n9288# A8 a_182_n9288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1377 a_1898_n71342# a_1848_n66# a_1766_n71342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1378 word656 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1379 word947 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1380 GND A4 word15 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1381 GND A3 word343 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1382 word597 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1383 word892 A0 a_2294_n126864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1384 word936 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1385 GND A2 word1008 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1386 word9 a_2376_n66# a_2294_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1387 a_1634_n17808# a_1584_n66# a_1370_n17808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1388 word877 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1389 a_578_n66372# a_528_n66# a_314_n66372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1390 word658 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1391 a_182_n10140# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1392 a_50_n88666# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1393 a_50_n97044# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1394 a_578_n57994# a_528_n66# a_314_n57994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1395 a_1238_n47912# A5 a_842_n47912# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1396 a_842_n67650# a_792_n66# a_578_n67650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1397 word165 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1398 word224 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1399 a_1898_n31440# a_1848_n66# a_1634_n31440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1400 GND A0 word344 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1401 a_50_n123598# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1402 word375 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1403 GND A0 word502 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1404 word556 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1405 a_314_n141206# a_264_n66# a_50_n141206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1406 a_1106_n144614# a_1056_n66# a_842_n144614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1407 a_314_n132828# a_264_n66# a_50_n132828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1408 word368 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1409 word653 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1410 word908 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1411 word221 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1412 a_842_n106558# a_792_n66# a_578_n106558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1413 a_578_n26470# a_528_n66# a_446_n26470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1414 GND A3 word177 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1415 word429 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1416 a_974_n74040# A6 a_710_n74040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1417 word726 A0 a_2162_n103292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1418 a_182_n56574# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1419 GND A3 word118 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1420 a_1502_n38682# A4 a_1238_n38682# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1421 a_314_n109966# a_264_n66# a_50_n109966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1422 a_314_n118344# a_264_n66# a_50_n118344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1423 GND A6 word549 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1424 a_1898_n86252# a_1848_n66# a_1634_n86252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1425 a_710_n12412# A7 a_446_n12412# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1426 a_578_n95766# a_528_n66# a_446_n95766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1427 word711 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1428 GND A2 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1429 word702 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1430 a_842_n35700# a_792_n66# a_578_n35700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1431 word268 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1432 word844 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1433 a_1634_n63532# a_1584_n66# a_1370_n63532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1434 word531 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1435 word982 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1436 a_182_n25050# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1437 GND A4 word544 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1438 word1007 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1439 word172 A0 a_2294_n24624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1440 word150 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1441 a_314_n54586# a_264_n66# a_182_n54586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1442 word830 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1443 a_1634_n113232# a_1584_n66# a_1370_n113232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1444 a_1898_n46350# a_1848_n66# a_1766_n46350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1445 word428 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1446 a_842_n144330# a_792_n66# a_578_n144330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1447 word35 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1448 word992 A0 a_2294_n141064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1449 GND A6 word781 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1450 word101 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1451 GND A3 word384 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1452 word638 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1453 word110 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1454 a_974_n110108# A6 a_710_n110108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1455 word760 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1456 word473 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1457 a_974_n42090# A6 a_710_n42090# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1458 word414 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1459 a_710_n41806# A7 a_314_n41806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1460 word918 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1461 word15 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1462 a_578_n72194# a_528_n66# a_314_n72194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1463 GND A5 word322 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1464 a_50_n94488# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1465 word534 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1466 a_2162_n14826# a_2112_n66# a_1898_n14826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1467 a_2162_n23204# a_2112_n66# a_2030_n23204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1468 a_1634_n92926# a_1584_n66# a_1502_n92926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1469 GND A2 word888 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1470 word816 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1471 word757 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1472 a_1634_n31582# a_1584_n66# a_1370_n31582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1473 word538 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1474 word315 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1475 word374 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1476 a_1634_n142626# a_1584_n66# a_1502_n142626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1477 word367 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1478 a_1898_n14400# a_1848_n66# a_1766_n14400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1479 a_1238_n22210# A5 a_974_n22210# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1480 word308 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1481 a_314_n69496# a_264_n66# a_182_n69496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1482 GND A9 word93 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1483 a_182_n62396# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1484 a_2294_n21216# A1 a_1898_n21216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1485 a_314_n115788# a_264_n66# a_50_n115788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1486 a_314_n124166# a_264_n66# a_50_n124166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1487 a_1634_n119764# a_1584_n66# a_1502_n119764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1488 a_2294_n12838# A1 a_2030_n12838# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1489 a_1898_n92074# a_1848_n66# a_1766_n92074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1490 word371 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1491 GND A3 word548 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1492 a_1898_n83696# a_1848_n66# a_1634_n83696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1493 a_1238_n91506# A5 a_974_n91506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1494 GND A5 word156 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1495 a_1766_n128426# A3 a_1502_n128426# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1496 GND A6 word827 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1497 a_1238_n21784# A5 a_974_n21784# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1498 a_1238_n30162# A5 a_842_n30162# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1499 a_2294_n90512# A1 a_1898_n90512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1500 a_974_n116640# A6 a_710_n116640# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1501 a_1634_n38540# a_1584_n66# a_1502_n38540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1502 word309 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1503 a_2030_n47202# A2 a_1634_n47202# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1504 word1023 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1505 a_2030_n38824# A2 a_1766_n38824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1506 a_2162_n123314# a_2112_n66# a_2030_n123314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1507 a_1634_n60976# a_1584_n66# a_1502_n60976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1508 a_1238_n77022# A5 a_974_n77022# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1509 GND A4 word585 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1510 a_2162_n38114# a_2112_n66# a_2030_n38114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1511 word741 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1512 a_1634_n110676# a_1584_n66# a_1502_n110676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1513 word90 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1514 word574 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1515 word411 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1516 word484 A0 a_2294_n68928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1517 GND A9 word31 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1518 word479 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1519 a_1502_n82276# A4 a_1238_n82276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1520 word210 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1521 a_1502_n73898# A4 a_1238_n73898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1522 GND A5 word205 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1523 a_446_n19512# A8 a_182_n19512# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1524 a_1238_n37120# A5 a_974_n37120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1525 a_842_n127290# a_792_n66# a_710_n127290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1526 GND A3 word323 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1527 GND A9 word198 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1528 a_314_n139076# a_264_n66# a_50_n139076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1529 GND A9 word139 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1530 a_2294_n36126# A1 a_1898_n36126# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1531 word639 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1532 word697 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1533 GND A9 word356 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1534 a_2030_n136946# A2 a_1766_n136946# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1535 word46 A0 a_2162_n6732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1536 word189 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1537 a_2030_n15252# A2 a_1634_n15252# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1538 GND A5 word261 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1539 word948 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1540 GND A5 word202 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1541 a_2162_n67508# a_2112_n66# a_2030_n67508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1542 a_1238_n36694# A5 a_974_n36694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1543 word677 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1544 a_446_n10424# A8 a_182_n10424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1545 word318 A0 a_2162_n45356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1546 word727 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1547 GND A9 word75 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1548 word254 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1549 a_1106_n133396# a_1056_n66# a_974_n133396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1550 word195 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1551 word679 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1552 word67 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1553 word247 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1554 GND A3 word530 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1555 GND A9 word405 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1556 word188 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1557 a_2294_n65520# A1 a_1898_n65520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1558 a_1502_n97186# A4 a_1106_n97186# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1559 GND A1 word729 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1560 a_1766_n134248# A3 a_1370_n134248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1561 a_1238_n101304# A5 a_842_n101304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1562 a_1766_n125870# A3 a_1370_n125870# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1563 GND A2 word96 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1564 a_2030_n44646# A2 a_1634_n44646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1565 a_578_n106842# a_528_n66# a_446_n106842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1566 a_2030_n104996# A2 a_1766_n104996# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1567 GND A5 word468 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1568 GND A5 word527 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1569 word431 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1570 a_1238_n74466# A5 a_974_n74466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1571 word870 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1572 a_3292_164# A1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X1573 word723 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1574 GND A9 word461 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1575 a_710_n115504# A7 a_314_n115504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1576 a_1502_n118912# A4 a_1238_n118912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1577 a_1766_n30304# A3 a_1370_n30304# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1578 a_710_n48054# A7 a_314_n48054# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1579 GND A8 word41 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1580 a_2294_n73472# A1 a_1898_n73472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1581 a_710_n39676# A7 a_314_n39676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1582 word584 A0 a_2294_n83128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1583 a_2162_n106274# a_2112_n66# a_2030_n106274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1584 word993 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1585 a_1634_n99174# a_1584_n66# a_1370_n99174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1586 a_446_n16956# A8 a_182_n16956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1587 a_446_n25334# A8 a_182_n25334# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1588 GND A1 word136 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1589 GND A7 word770 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1590 GND A8 word631 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1591 GND A9 word239 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1592 GND A2 word362 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1593 GND A9 word180 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1594 a_2030_n82418# A2 a_1766_n82418# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1595 word773 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1596 a_578_n144614# a_528_n66# a_314_n144614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1597 a_2030_n12696# A2 a_1634_n12696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1598 a_2030_n21074# A2 a_1766_n21074# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1599 word989 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1600 GND A8 word79 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1601 a_2162_n73330# a_2112_n66# a_2030_n73330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1602 GND A6 word914 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1603 GND A1 word893 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1604 word704 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1605 a_446_n104428# A8 a_50_n104428# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1606 GND A7 word826 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1607 GND A3 word996 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1608 a_1106_n6874# a_1056_n66# a_974_n6874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1609 a_2294_n19086# A1 a_1898_n19086# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1610 GND A2 word201 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1611 a_710_n77448# A7 a_446_n77448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1612 a_2030_n59556# A2 a_1766_n59556# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1613 word578 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1614 GND A1 word72 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1615 GND A6 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1616 word536 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1617 a_1634_n90086# a_1584_n66# a_1370_n90086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1618 word659 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1619 word975 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1620 word477 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1621 a_2030_n81992# A2 a_1766_n81992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1622 GND A8 word567 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1623 a_2162_n135668# a_2112_n66# a_2030_n135668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1624 word300 A0 a_2294_n42800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1625 GND A7 word262 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1626 word295 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1627 a_2294_n88382# A1 a_1898_n88382# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1628 word709 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1629 word27 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1630 a_1766_n36836# A3 a_1502_n36836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1631 GND A8 word76 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1632 a_2162_n81282# a_2112_n66# a_2030_n81282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1633 a_2294_n101446# A1 a_2030_n101446# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1634 word288 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1635 word557 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1636 word630 A0 a_2162_n89660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1637 a_1106_n17808# a_1056_n66# a_842_n17808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1638 GND A3 word774 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1639 a_2294_n139928# A1 a_2030_n139928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1640 a_2030_n50468# A2 a_1766_n50468# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1641 word715 a_2376_n66# a_2162_n101730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1642 word255 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1643 word559 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1644 GND A1 word68 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1645 GND A9 word344 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1646 GND A2 word467 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1647 GND A9 word502 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1648 a_1502_n133112# A4 a_1106_n133112# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1649 GND A4 word898 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1650 a_2162_n41380# a_2112_n66# a_2030_n41380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1651 a_2294_n48480# A1 a_1898_n48480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1652 a_2030_n88950# A2 a_1766_n88950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1653 a_710_n112948# A7 a_314_n112948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1654 a_1502_n124734# A4 a_1106_n124734# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1655 a_710_n121326# A7 a_314_n121326# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1656 GND A8 word23 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1657 a_710_n45498# A7 a_314_n45498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1658 a_1370_n35416# a_1320_n66# a_1106_n35416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1659 GND A8 word125 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1660 GND A8 word184 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1661 word750 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1662 word241 a_2376_n66# a_2294_n34422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1663 word252 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1664 a_2294_n130840# A1 a_2030_n130840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1665 a_446_n22778# A8 a_182_n22778# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1666 a_446_n31156# A8 a_182_n31156# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1667 GND A1 word177 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1668 word495 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1669 GND A6 word54 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1670 word464 A0 a_2294_n66088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1671 GND A8 word672 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1672 word873 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1673 a_446_n78016# A8 a_50_n78016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1674 GND A8 word742 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1675 GND A7 word42 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1676 GND A2 word674 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1677 word803 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1678 a_1238_n122036# A5 a_842_n122036# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1679 GND A3 word820 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1680 a_1106_n63532# a_1056_n66# a_974_n63532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1681 GND A9 word119 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1682 word879 a_2376_n66# a_2162_n125018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1683 a_1238_n113658# A5 a_974_n113658# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1684 GND A2 word242 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1685 a_2030_n65378# A2 a_1634_n65378# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1686 a_710_n83270# A7 a_446_n83270# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1687 a_1502_n101162# A4 a_1238_n101162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1688 a_578_n127574# a_528_n66# a_314_n127574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1689 a_2030_n57000# A2 a_1766_n57000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1690 word784 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1691 a_1238_n95198# A5 a_974_n95198# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1692 a_2162_n141490# a_2112_n66# a_2030_n141490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1693 GND A5 word906 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1694 a_1370_n122320# a_1320_n66# a_1238_n122320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1695 GND A7 word303 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1696 a_974_n5028# A6 a_710_n5028# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1697 a_50_n112806# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1698 a_1766_n51036# A3 a_1502_n51036# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1699 GND A1 word384 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1700 a_2162_n56290# a_2112_n66# a_2030_n56290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1701 GND A8 word69 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1702 word9 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1703 GND A0 word984 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1704 a_1106_n23630# a_1056_n66# a_974_n23630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1705 a_1106_n32008# a_1056_n66# a_842_n32008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1706 a_1370_n72762# a_1320_n66# a_1106_n72762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1707 GND A6 word143 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1708 a_1766_n89518# A3 a_1370_n89518# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1709 word937 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1710 a_1370_n130272# a_1320_n66# a_1238_n130272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1711 word878 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1712 a_1370_n121894# a_1320_n66# a_1238_n121894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1713 a_1766_n28174# A3 a_1502_n28174# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1714 word1010 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1715 GND A9 word57 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1716 GND A2 word449 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1717 GND A4 word939 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1718 GND A0 word920 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1719 GND A8 word225 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1720 word908 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1721 GND A1 word980 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1722 a_1238_n128568# A5 a_974_n128568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1723 GND A2 word347 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1724 a_974_n62822# A6 a_578_n62822# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1725 a_1106_n78442# a_1056_n66# a_974_n78442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1726 a_1766_n80430# A3 a_1370_n80430# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1727 GND A4 word837 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1728 word223 a_2376_n66# a_2162_n31866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1729 GND A7 word78 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1730 a_1370_n79720# a_1320_n66# a_1106_n79720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1731 word931 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1732 word682 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1733 GND A8 word555 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1734 word889 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1735 word623 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1736 GND A0 word818 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1737 GND A7 word349 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1738 GND A1 word548 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1739 word553 a_2376_n66# a_2294_n78726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1740 a_446_n4318# A8 a_182_n4318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1741 a_50_n127716# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1742 word121 a_2376_n66# a_2294_n17382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1743 a_446_n75460# A8 a_50_n75460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1744 a_1766_n57568# A3 a_1370_n57568# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1745 GND A1 word489 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1746 GND A7 word566 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1747 a_2294_n113800# A1 a_2030_n113800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1748 a_182_n13832# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1749 a_974_n22920# A6 a_578_n22920# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1750 word844 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1751 GND A8 word552 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1752 a_1106_n60976# a_1056_n66# a_974_n60976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1753 word785 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1754 a_1370_n145182# a_1320_n66# a_1106_n145182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1755 a_578_n61402# a_528_n66# a_314_n61402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1756 GND A2 word283 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1757 GND A4 word714 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1758 word751 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1759 a_578_n133396# a_528_n66# a_314_n133396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1760 a_446_n3892# A8 a_182_n3892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1761 GND A2 word554 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1762 GND A1 word425 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1763 GND A7 word285 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1764 word46 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1765 word457 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1766 a_974_n77732# A6 a_710_n77732# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1767 GND A7 word615 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1768 a_842_n70632# a_792_n66# a_578_n70632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1769 word387 a_2376_n66# a_2162_n55154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1770 a_50_n104144# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1771 word179 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1772 GND A0 word306 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1773 a_710_n119196# A7 a_314_n119196# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1774 a_182_n51604# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1775 a_314_n58704# a_264_n66# a_182_n58704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1776 a_1502_n33712# A4 a_1106_n33712# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1777 GND A1 word264 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1778 GND A5 word725 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1779 word667 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1780 a_2294_n137088# A1 a_1898_n137088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1781 word962 A0 a_2162_n136804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1782 a_182_n28742# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1783 GND A5 word19 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1784 a_842_n30730# a_792_n66# a_578_n30730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1785 word174 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1786 a_974_n37830# A6 a_710_n37830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1787 word890 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1788 GND A0 word84 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1789 word755 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1790 a_710_n9146# A7 a_446_n9146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1791 a_578_n67934# a_528_n66# a_314_n67934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1792 a_50_n98606# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1793 GND A3 word51 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1794 GND A4 word77 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1795 word61 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1796 word664 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1797 a_842_n16246# a_792_n66# a_710_n16246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1798 GND A0 word572 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1799 GND A0 word800 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1800 GND A7 a_528_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X1801 a_50_n133538# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1802 word811 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1803 a_1370_n93494# a_1320_n66# a_1238_n93494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1804 word752 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1805 GND A6 word289 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1806 a_842_n85542# a_792_n66# a_710_n85542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1807 a_578_n36410# a_528_n66# a_446_n36410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1808 a_50_n119054# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1809 word851 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1810 a_1898_n40954# a_1848_n66# a_1634_n40954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1811 word501 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1812 word796 A0 a_2294_n113232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1813 a_182_n66514# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1814 word442 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1815 a_314_n119906# a_264_n66# a_50_n119906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1816 GND A6 word560 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1817 GND A5 word988 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1818 word277 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1819 a_1634_n2330# a_1584_n66# a_1502_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1820 a_2294_n3750# A1 a_2030_n3750# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1821 GND A2 word595 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1822 word781 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1823 GND A6 word128 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1824 word562 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1825 word722 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1826 GND A2 word794 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1827 a_578_n35984# a_528_n66# a_446_n35984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1828 a_50_n75034# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1829 a_842_n54018# a_792_n66# a_710_n54018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1830 a_842_n45640# a_792_n66# a_710_n45640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1831 word279 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1832 a_1106_n99174# a_1056_n66# a_974_n99174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1833 word855 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1834 GND A0 word130 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1835 word369 a_2376_n66# a_2294_n52598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1836 a_182_n8436# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1837 a_50_n101588# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1838 word220 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1839 word1018 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1840 a_314_n64526# a_264_n66# a_182_n64526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1841 a_314_n110818# a_264_n66# a_50_n110818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1842 word699 a_2376_n66# a_2162_n99458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1843 word498 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1844 GND A0 word964 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1845 a_842_n53592# a_792_n66# a_710_n53592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1846 a_1766_n78300# A3 a_1502_n78300# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1847 GND A0 word618 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1848 a_182_n34564# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1849 GND A4 word611 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1850 word484 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1851 a_1370_n9004# a_1320_n66# a_1106_n9004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1852 word215 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1853 GND A6 word394 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1854 a_1106_n90086# a_1056_n66# a_842_n90086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1855 word396 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1856 word606 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1857 a_710_n6590# A7 a_446_n6590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1858 GND A4 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1859 word842 A0 a_2162_n119764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1860 GND A3 word33 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1861 a_842_n13690# a_792_n66# a_710_n13690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1862 word236 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1863 word635 a_2376_n66# a_2162_n90370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1864 word886 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1865 word827 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1866 GND A2 word899 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1867 word608 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1868 a_578_n59272# a_528_n66# a_314_n59272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1869 GND A4 word389 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1870 a_974_n98464# A6 a_578_n98464# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1871 a_842_n122320# a_792_n66# a_710_n122320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1872 a_842_n82986# a_792_n66# a_710_n82986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1873 a_50_n116498# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1874 GND A0 word452 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1875 a_182_n63958# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1876 a_182_n72336# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1877 GND A3 word229 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1878 a_314_n134106# a_264_n66# a_50_n134106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1879 word662 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1880 word778 A0 a_2162_n110676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1881 a_314_n125728# a_264_n66# a_50_n125728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1882 word318 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1883 word259 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1884 a_974_n20080# A6 a_578_n20080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1885 a_578_n19370# a_528_n66# a_446_n19370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1886 a_1502_n5738# A4 a_1106_n5738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1887 GND A6 word169 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1888 word171 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1889 a_1238_n40102# A5 a_974_n40102# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1890 a_842_n121894# a_792_n66# a_710_n121894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1891 a_182_n49474# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1892 a_1238_n31724# A5 a_842_n31724# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1893 a_974_n80998# A6 a_710_n80998# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1894 a_578_n97044# a_528_n66# a_446_n97044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1895 a_1898_n79152# a_1848_n66# a_1634_n79152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1896 GND A4 word655 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1897 GND A6 word657 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1898 a_182_n5880# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1899 word151 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1900 a_314_n61970# a_264_n66# a_182_n61970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1901 a_314_n70348# a_264_n66# a_182_n70348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1902 GND A4 word164 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1903 a_974_n134532# A6 a_578_n134532# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1904 a_842_n28600# a_792_n66# a_578_n28600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1905 word481 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1906 word341 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1907 word735 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1908 a_1634_n56432# a_1584_n66# a_1502_n56432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1909 a_1502_n92216# A4 a_1238_n92216# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1910 word60 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1911 word122 A0 a_2162_n17524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1912 a_1502_n83838# A4 a_1238_n83838# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1913 word957 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1914 a_182_n40386# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1915 a_314_n47486# a_264_n66# a_182_n47486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1916 GND A4 word652 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1917 a_1634_n106132# a_1584_n66# a_1502_n106132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1918 GND A2 word16 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1919 a_1106_n105564# a_1056_n66# a_842_n105564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1920 word437 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1921 a_842_n137230# a_792_n66# a_578_n137230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1922 a_1898_n70064# a_1848_n66# a_1634_n70064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1923 word938 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1924 a_1502_n69354# A4 a_1106_n69354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1925 word546 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1926 word95 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1927 GND A5 word331 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1928 word868 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1929 GND A5 word272 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1930 word649 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1931 a_842_n145182# a_792_n66# a_578_n145182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1932 a_578_n65094# a_528_n66# a_314_n65094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1933 a_1238_n46634# A5 a_842_n46634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1934 a_1238_n55012# A5 a_974_n55012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1935 GND A4 word430 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1936 word590 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1937 a_50_n87388# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1938 word116 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1939 word583 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1940 a_1634_n85826# a_1584_n66# a_1370_n85826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1941 GND A2 word65 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1942 a_1634_n24482# a_1584_n66# a_1502_n24482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1943 GND A4 word269 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1944 a_1502_n51888# A4 a_1106_n51888# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1945 a_1502_n60266# A4 a_1106_n60266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1946 a_314_n131550# a_264_n66# a_50_n131550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1947 a_1106_n143336# a_1056_n66# a_842_n143336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1948 a_1634_n135526# a_1584_n66# a_1370_n135526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1949 a_1106_n134958# a_1056_n66# a_974_n134958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1950 word644 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1951 word359 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1952 word300 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1953 a_1898_n114652# a_1848_n66# a_1766_n114652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1954 word317 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1955 a_842_n105280# a_792_n66# a_578_n105280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1956 GND A7 word791 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1957 a_182_n55296# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1958 a_314_n117066# a_264_n66# a_50_n117066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1959 a_2030_n123314# A2 a_1766_n123314# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1960 word483 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1961 a_2030_n114936# A2 a_1634_n114936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1962 a_710_n11134# A7 a_446_n11134# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1963 a_578_n94488# a_528_n66# a_446_n94488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1964 a_1238_n84406# A5 a_842_n84406# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1965 GND A3 word597 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1966 GND A3 word656 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1967 a_974_n109540# A6 a_710_n109540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1968 a_1766_n143762# A3 a_1370_n143762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1969 a_710_n49616# A7 a_314_n49616# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1970 word382 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1971 word973 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1972 a_974_n131976# A6 a_578_n131976# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1973 a_1634_n53876# a_1584_n66# a_1370_n53876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1974 word463 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1975 word914 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1976 word695 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1977 a_2162_n107836# a_2112_n66# a_1898_n107836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1978 word996 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1979 word104 A0 a_2294_n14968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1980 word99 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1981 a_1634_n103576# a_1584_n66# a_1370_n103576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1982 a_974_n117492# A6 a_710_n117492# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1983 GND A3 word375 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1984 a_2294_n43510# A1 a_2030_n43510# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1985 word464 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1986 word843 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1987 a_1766_n112238# A3 a_1370_n112238# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1988 word587 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1989 a_1898_n129562# a_1848_n66# a_1634_n129562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1990 a_710_n40528# A7 a_314_n40528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1991 a_2030_n31014# A2 a_1634_n31014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1992 word850 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1993 word715 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1994 word589 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1995 GND A9 word306 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X1996 a_2030_n129846# A2 a_1766_n129846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1997 a_2162_n13548# a_2112_n66# a_1898_n13548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X1998 a_2294_n51462# A1 a_2030_n51462# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X1999 a_710_n17666# A7 a_446_n17666# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2000 word297 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2001 word370 A0 a_2162_n52740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2002 word898 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2003 word779 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2004 a_1238_n29594# A5 a_842_n29594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2005 GND A8 word146 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2006 a_2162_n82844# a_2112_n66# a_1898_n82844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2007 a_2294_n89944# A1 a_2030_n89944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2008 word487 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2009 word358 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2010 a_1634_n77164# a_1584_n66# a_1370_n77164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2011 word627 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2012 a_1898_n120474# a_1848_n66# a_1634_n120474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2013 word299 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2014 a_710_n86962# A7 a_446_n86962# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2015 GND A6 word920 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2016 word268 A0 a_2294_n38256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2017 GND A9 word84 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2018 GND A3 word150 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2019 a_1106_n126296# a_1056_n66# a_842_n126296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2020 a_2294_n11560# A1 a_2030_n11560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2021 a_2030_n60408# A2 a_1634_n60408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2022 word426 A0 a_2162_n60692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2023 GND A5 word579 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2024 word629 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2025 a_2030_n120758# A2 a_1766_n120758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2026 GND A5 word147 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2027 GND A3 word480 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2028 GND A6 word818 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2029 GND A5 word88 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2030 a_1766_n118770# A3 a_1502_n118770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2031 a_2294_n80856# A1 a_2030_n80856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2032 a_2030_n106274# A2 a_1634_n106274# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2033 word364 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2034 word563 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2035 word1014 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2036 word381 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2037 word879 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2038 a_2162_n122036# a_2112_n66# a_2030_n122036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2039 a_1238_n58988# A5 a_974_n58988# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2040 a_1238_n67366# A5 a_842_n67366# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2041 GND A5 word576 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2042 word732 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2043 a_2162_n113658# a_2112_n66# a_1898_n113658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2044 GND A9 word411 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2045 a_1766_n23204# A3 a_1502_n23204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2046 a_2162_n28458# a_2112_n66# a_1898_n28458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2047 word565 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2048 a_446_n32718# A8 a_182_n32718# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2049 a_1766_n14826# A3 a_1502_n14826# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2050 word534 A0 a_2162_n76028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2051 GND A9 word22 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2052 word943 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2053 word876 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2054 GND A8 word251 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2055 a_2162_n97754# a_2112_n66# a_1898_n97754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2056 a_2294_n117918# A1 a_1898_n117918# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2057 a_446_n18234# A8 a_182_n18234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2058 GND A1 a_2112_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X2059 GND A7 word53 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2060 GND A7 word878 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2061 GND A9 word189 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2062 GND A2 word312 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2063 a_2030_n75318# A2 a_1766_n75318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2064 GND A9 word130 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2065 a_2030_n135668# A2 a_1634_n135668# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2066 a_578_n137514# a_528_n66# a_314_n137514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2067 a_1502_n111102# A4 a_1238_n111102# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2068 GND A4 word743 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2069 a_2294_n26470# A1 a_2030_n26470# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2070 a_1370_n13406# a_1320_n66# a_1238_n13406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2071 word939 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2072 word156 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2073 a_1106_n8152# a_1056_n66# a_974_n8152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2074 a_2294_n95766# A1 a_2030_n95766# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2075 GND A1 word1001 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2076 GND A3 word946 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2077 word469 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2078 word609 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2079 GND A3 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2080 GND A8 word517 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2081 word250 A0 a_2162_n35700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2082 a_1370_n140212# a_1320_n66# a_1238_n140212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2083 a_1370_n131834# a_1320_n66# a_1238_n131834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2084 a_1766_n29736# A3 a_1370_n29736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2085 GND A9 word68 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2086 GND A1 word720 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2087 GND A3 word724 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2088 GND A6 word800 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2089 a_1106_n41522# a_1056_n66# a_974_n41522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2090 word205 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2091 a_2030_n43368# A2 a_1766_n43368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2092 a_578_n105564# a_528_n66# a_446_n105564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2093 a_1370_n108972# a_1320_n66# a_1106_n108972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2094 GND A5 word400 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2095 GND A5 word459 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2096 word363 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2097 GND A2 word417 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2098 a_1238_n73188# A5 a_974_n73188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2099 a_1238_n138508# A5 a_842_n138508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2100 word293 a_2376_n66# a_2294_n41806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2101 a_710_n114226# A7 a_314_n114226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2102 word714 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2103 GND A9 word452 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2104 GND A1 word229 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2105 GND A7 word89 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2106 GND A1 word776 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2107 a_710_n38398# A7 a_314_n38398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2108 a_1766_n20648# A3 a_1370_n20648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2109 GND A3 word721 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2110 GND A8 word134 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2111 word721 a_2376_n66# a_2294_n102582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2112 word202 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2113 GND A7 word636 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2114 word925 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2115 word191 a_2376_n66# a_2162_n27322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2116 a_2294_n132118# A1 a_2030_n132118# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2117 word782 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2118 a_446_n24056# A8 a_182_n24056# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2119 a_446_n15678# A8 a_182_n15678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2120 GND A1 word13 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2121 GND A6 word63 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2122 word445 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2123 word855 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2124 GND A8 word622 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2125 word956 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2126 GND A2 word353 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2127 a_1106_n70916# a_1056_n66# a_842_n70916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2128 a_2030_n81140# A2 a_1634_n81140# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2129 a_2030_n141490# A2 a_1766_n141490# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2130 word823 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2131 a_578_n143336# a_528_n66# a_314_n143336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2132 a_2162_n89092# a_2112_n66# a_2030_n89092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2133 a_578_n134958# a_528_n66# a_314_n134958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2134 a_2294_n109256# A1 a_2030_n109256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2135 word53 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2136 a_446_n84974# A8 a_50_n84974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2137 a_446_n93352# A8 a_50_n93352# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2138 GND A2 word624 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2139 GND A8 word70 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2140 GND A7 word355 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2141 a_446_n103150# A8 a_50_n103150# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2142 GND A1 word825 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2143 GND A3 word770 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2144 a_974_n40812# A6 a_710_n40812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2145 GND A2 word192 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2146 a_710_n76170# A7 a_446_n76170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2147 GND A3 word928 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2148 a_1106_n5596# a_1056_n66# a_974_n5596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2149 a_1370_n57710# a_1320_n66# a_1238_n57710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2150 a_2030_n58278# A2 a_1634_n58278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2151 word987 a_2376_n66# a_2162_n140354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2152 word527 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2153 word734 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2154 GND A1 word393 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2155 word989 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2156 a_50_n105706# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2157 a_2294_n100168# A1 a_2030_n100168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2158 a_1106_n16530# a_1056_n66# a_842_n16530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2159 word828 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2160 word550 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2161 GND A2 word458 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2162 word960 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2163 GND A5 word851 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2164 GND A5 word792 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2165 a_2030_n96050# A2 a_1766_n96050# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2166 a_1502_n123456# A4 a_1106_n123456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2167 a_710_n120048# A7 a_314_n120048# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2168 a_1106_n24482# a_1056_n66# a_974_n24482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2169 a_710_n111670# A7 a_314_n111670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2170 GND A8 word14 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2171 a_446_n99884# A8 a_50_n99884# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2172 a_1370_n25760# a_1320_n66# a_1106_n25760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2173 GND A8 word175 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2174 GND A0 word870 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2175 a_842_n17808# a_792_n66# a_710_n17808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2176 word302 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2177 a_974_n55722# A6 a_578_n55722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2178 word173 a_2376_n66# a_2294_n24766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2179 a_1766_n73330# A3 a_1502_n73330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2180 word1016 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2181 word881 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2182 GND A1 word168 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2183 word822 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2184 a_446_n21500# A8 a_182_n21500# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2185 GND A1 word109 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2186 GND A6 word45 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2187 GND A8 word663 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2188 GND A8 word604 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2189 GND A0 word768 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2190 GND A8 word733 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2191 GND A0 word926 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2192 word862 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2193 a_710_n1620# A7 a_446_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2194 GND A1 word656 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2195 GND A7 word516 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2196 a_2294_n115078# A1 a_2030_n115078# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2197 a_578_n140780# a_528_n66# a_314_n140780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2198 a_446_n90796# A8 a_50_n90796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2199 GND A1 word597 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2200 a_2294_n768# A1 a_1898_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2201 GND A2 word665 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2202 a_1106_n62254# a_1056_n66# a_974_n62254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2203 GND A9 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2204 a_1238_n112380# A5 a_974_n112380# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2205 a_446_n484# A8 a_182_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2206 GND A2 word233 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2207 GND A6 word139 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2208 a_1106_n53876# a_1056_n66# a_842_n53876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2209 a_2030_n64100# A2 a_1766_n64100# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2210 word509 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2211 word439 a_2376_n66# a_2162_n62538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2212 GND A0 word704 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2213 GND A6 word686 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2214 GND A5 word897 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2215 a_50_n111528# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2216 a_1502_n138366# A4 a_1238_n138366# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2217 a_710_n126580# A7 a_314_n126580# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2218 GND A2 word762 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2219 a_974_n23772# A6 a_578_n23772# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2220 a_1766_n41380# A3 a_1502_n41380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2221 a_2162_n1194# a_2112_n66# a_1898_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2222 GND A4 word193 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2223 a_1370_n49048# a_1320_n66# a_1238_n49048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2224 a_1370_n71484# a_1320_n66# a_1106_n71484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2225 word337 a_2376_n66# a_2294_n48054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2226 GND A0 word256 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2227 GND A4 word681 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2228 a_182_n44504# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2229 word287 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2230 GND A2 word499 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2231 GND A6 word405 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2232 word967 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2233 GND A2 word440 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2234 a_1898_n65804# a_1848_n66# a_1634_n65804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2235 GND A7 word621 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2236 GND A4 word930 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2237 a_1766_n96192# A3 a_1502_n96192# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2238 word912 A0 a_2294_n129704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2239 a_578_n22352# a_528_n66# a_446_n22352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2240 GND A5 word28 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2241 a_842_n32008# a_792_n66# a_578_n32008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2242 word124 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2243 a_974_n39108# A6 a_710_n39108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2244 word29 a_2376_n66# a_2294_n4318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2245 a_974_n61544# A6 a_578_n61544# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2246 word840 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2247 a_578_n69212# a_528_n66# a_314_n69212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2248 GND A2 word338 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2249 a_1106_n68786# a_1056_n66# a_842_n68786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2250 GND A4 word769 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2251 a_314_n42516# a_264_n66# a_182_n42516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2252 word880 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2253 GND A4 word32 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2254 a_1370_n17098# a_1320_n66# a_1106_n17098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2255 GND A0 word750 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2256 GND A8 word645 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2257 a_446_n3040# A8 a_182_n3040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2258 a_50_n126438# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2259 a_1898_n8720# a_1848_n66# a_1634_n8720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2260 GND A7 word340 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2261 GND A0 word522 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2262 a_842_n31582# a_792_n66# a_578_n31582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2263 a_974_n38682# A6 a_710_n38682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2264 GND A1 word480 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2265 word848 A0 a_2294_n120616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2266 a_1766_n2472# A3 a_1370_n2472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2267 word761 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2268 a_182_n12554# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2269 GND A4 word456 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2270 a_1370_n86394# a_1320_n66# a_1238_n86394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2271 word329 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2272 a_578_n29310# a_528_n66# a_446_n29310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2273 GND A0 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2274 GND A6 word180 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2275 word241 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2276 a_578_n60124# a_528_n66# a_314_n60124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2277 word742 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2278 a_842_n140212# a_792_n66# a_578_n140212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2279 a_182_n59414# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2280 a_50_n82418# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2281 a_1898_n33854# a_1848_n66# a_1634_n33854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2282 word746 A0 a_2162_n106132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2283 word81 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2284 a_578_n98606# a_528_n66# a_446_n98606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2285 GND A2 word545 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2286 GND A2 word744 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2287 word731 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2288 GND A2 word803 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2289 a_578_n28884# a_528_n66# a_446_n28884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2290 a_314_n71910# a_264_n66# a_182_n71910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2291 a_1238_n18802# A5 a_974_n18802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2292 GND A4 word234 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2293 a_842_n108972# a_792_n66# a_578_n108972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2294 a_50_n81992# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2295 a_1766_n9430# A3 a_1502_n9430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2296 a_974_n76454# A6 a_710_n76454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2297 word446 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2298 a_842_n100310# a_792_n66# a_578_n100310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2299 word805 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2300 word319 a_2376_n66# a_2162_n45498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2301 a_314_n57426# a_264_n66# a_182_n57426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2302 GND A0 word238 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2303 a_182_n41948# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2304 a_182_n50326# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2305 a_1502_n32434# A4 a_1106_n32434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2306 a_1106_n115504# a_1056_n66# a_974_n115504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2307 word448 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2308 word55 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2309 a_842_n46492# a_792_n66# a_710_n46492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2310 word286 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2311 a_1898_n71626# a_1848_n66# a_1766_n71626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2312 a_1238_n1762# A5 a_974_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2313 word658 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2314 word861 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2315 a_1898_n10282# a_1848_n66# a_1766_n10282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2316 a_182_n27464# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2317 word165 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2318 GND A2 word1010 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2319 a_578_n66656# a_528_n66# a_314_n66656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2320 word660 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2321 a_50_n97328# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2322 a_1898_n48764# a_1848_n66# a_1766_n48764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2323 a_50_n88950# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2324 word52 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2325 word585 a_2376_n66# a_2294_n83270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2326 word653 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2327 a_974_n112522# A6 a_710_n112522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2328 a_50_n132260# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2329 word221 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2330 a_1502_n70206# A4 a_1106_n70206# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2331 GND A0 word504 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2332 word558 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2333 word429 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2334 word802 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2335 word370 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2336 word910 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2337 a_842_n84264# a_792_n66# a_710_n84264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2338 word551 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2339 a_50_n109398# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2340 word275 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2341 GND A0 word402 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2342 word223 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2343 word783 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2344 a_182_n65236# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2345 GND A3 word179 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2346 a_1502_n47344# A4 a_1238_n47344# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2347 a_314_n127006# a_264_n66# a_50_n127006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2348 a_182_n56858# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2349 word433 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2350 a_314_n118628# a_264_n66# a_50_n118628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2351 word728 A0 a_2294_n103576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2352 word268 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2353 word391 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2354 word713 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2355 word426 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2356 word966 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2357 GND A2 word785 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2358 a_842_n123172# a_792_n66# a_710_n123172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2359 word270 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2360 word428 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2361 a_974_n73898# A6 a_710_n73898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2362 word984 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2363 a_182_n7158# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2364 a_314_n63248# a_264_n66# a_182_n63248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2365 word101 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2366 word174 A0 a_2162_n24908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2367 word1009 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2368 a_314_n54870# a_264_n66# a_182_n54870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2369 a_1634_n113516# a_1584_n66# a_1370_n113516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2370 word110 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2371 a_974_n127432# A6 a_578_n127432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2372 word162 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2373 word326 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2374 a_1634_n49332# a_1584_n66# a_1370_n49332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2375 GND A0 word668 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2376 word990 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2377 a_2030_n5170# A2 a_1766_n5170# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2378 word103 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2379 word994 A0 a_2162_n141348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2380 word475 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2381 a_1898_n139502# a_1848_n66# a_1766_n139502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2382 a_182_n33286# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2383 a_1502_n15394# A4 a_1106_n15394# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2384 a_2030_n101304# A2 a_1634_n101304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2385 word387 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2386 word920 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2387 word166 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2388 a_578_n72478# a_528_n66# a_314_n72478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2389 a_1898_n54586# a_1848_n66# a_1634_n54586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2390 word538 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2391 GND A3 word501 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2392 GND A0 word56 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2393 word227 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2394 word367 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2395 word818 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2396 GND A2 word890 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2397 a_1634_n31866# a_1584_n66# a_1370_n31866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2398 a_1634_n40244# a_1584_n66# a_1370_n40244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2399 word540 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2400 word599 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2401 word759 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2402 a_842_n138082# a_792_n66# a_578_n138082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2403 a_1238_n39534# A5 a_974_n39534# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2404 a_1634_n142910# a_1584_n66# a_1502_n142910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2405 a_974_n97186# A6 a_578_n97186# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2406 a_1898_n130414# a_1848_n66# a_1766_n130414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2407 a_842_n90086# a_792_n66# a_710_n90086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2408 word533 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2409 a_1634_n78726# a_1584_n66# a_1502_n78726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2410 a_182_n71058# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2411 a_1634_n17382# a_1584_n66# a_1370_n17382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2412 a_1106_n136236# a_1056_n66# a_974_n136236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2413 a_182_n62680# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2414 a_314_n69780# a_264_n66# a_182_n69780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2415 word274 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2416 word496 A0 a_2294_n70632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2417 a_314_n124450# a_264_n66# a_50_n124450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2418 word309 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2419 a_2162_n69922# a_2112_n66# a_2030_n69922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2420 a_1898_n107552# a_1848_n66# a_1766_n107552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2421 GND A5 word217 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2422 a_1898_n83980# a_1848_n66# a_1634_n83980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2423 word1007 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2424 GND A5 word158 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2425 GND A6 word829 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2426 a_1238_n30446# A5 a_842_n30446# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2427 a_182_n48196# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2428 word493 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2429 GND A9 word151 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2430 a_2030_n116214# A2 a_1766_n116214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2431 word271 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2432 a_1238_n77306# A5 a_974_n77306# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2433 GND A5 word646 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2434 word743 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2435 GND A9 word481 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2436 word83 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2437 word210 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2438 a_2294_n76312# A1 a_2030_n76312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2439 GND A3 word547 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2440 a_2162_n60834# a_2112_n66# a_2030_n60834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2441 a_2294_n67934# A1 a_1898_n67934# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2442 word332 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2443 a_1766_n136662# A3 a_1502_n136662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2444 a_974_n133254# A6 a_578_n133254# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2445 a_1634_n110960# a_1584_n66# a_1502_n110960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2446 GND A0 word650 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2447 a_1634_n46776# a_1584_n66# a_1502_n46776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2448 word413 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2449 GND A4 word485 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2450 a_1502_n82560# A4 a_1238_n82560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2451 a_2162_n109114# a_2112_n66# a_1898_n109114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2452 a_1898_n145324# a_1848_n66# a_1634_n145324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2453 word639 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2454 a_2162_n37972# a_2112_n66# a_2030_n37972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2455 GND A3 word325 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2456 a_1502_n59698# A4 a_1106_n59698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2457 a_314_n139360# a_264_n66# a_50_n139360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2458 a_1766_n105138# A3 a_1502_n105138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2459 word699 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2460 GND A0 word38 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2461 a_1898_n98890# a_1848_n66# a_1766_n98890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2462 word859 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2463 word800 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2464 word724 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2465 GND A5 word263 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2466 a_2162_n100026# a_2112_n66# a_1898_n100026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2467 word640 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2468 a_1238_n36978# A5 a_974_n36978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2469 word598 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2470 GND A1 word1012 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2471 GND A9 word256 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2472 a_446_n10708# A8 a_182_n10708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2473 word679 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2474 a_2162_n138508# a_2112_n66# a_1898_n138508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2475 a_2294_n35984# A1 a_1898_n35984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2476 word107 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2477 word247 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2478 word320 A0 a_2294_n45640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2479 a_1106_n142058# a_1056_n66# a_842_n142058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2480 a_2162_n84122# a_2112_n66# a_1898_n84122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2481 word729 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2482 a_1106_n133680# a_1056_n66# a_974_n133680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2483 word721 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2484 GND A8 word96 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2485 a_1898_n113374# a_1848_n66# a_1634_n113374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2486 a_446_n106842# A8 a_50_n106842# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2487 GND A6 word929 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2488 word249 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2489 a_710_n79862# A7 a_446_n79862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2490 a_1502_n97470# A4 a_1106_n97470# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2491 GND A7 word782 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2492 a_2030_n122036# A2 a_1634_n122036# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2493 GND A3 word100 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2494 word376 A0 a_2294_n53592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2495 a_2030_n44930# A2 a_1634_n44930# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2496 GND A5 word470 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2497 GND A5 word529 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2498 a_1238_n83128# A5 a_842_n83128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2499 a_1238_n74750# A5 a_974_n74750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2500 GND A3 word647 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2501 GND A6 word768 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2502 a_2162_n44220# a_2112_n66# a_1898_n44220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2503 a_2294_n82134# A1 a_2030_n82134# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2504 GND A6 word926 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2505 GND A9 word463 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2506 a_710_n48338# A7 a_314_n48338# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2507 GND A8 word43 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2508 word373 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2509 GND A3 word791 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2510 a_710_n39960# A7 a_314_n39960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2511 word513 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2512 word964 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2513 a_974_n130698# A6 a_578_n130698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2514 word791 a_2376_n66# a_2162_n112522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2515 word331 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2516 a_2030_n52882# A2 a_1766_n52882# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2517 word154 A0 a_2162_n22068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2518 GND A5 word526 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2519 word987 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2520 a_1634_n102298# a_1584_n66# a_1502_n102298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2521 a_1898_n142768# a_1848_n66# a_1634_n142768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2522 word793 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2523 a_446_n25618# A8 a_182_n25618# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2524 a_1766_n16104# A3 a_1370_n16104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2525 a_2162_n52172# a_2112_n66# a_1898_n52172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2526 a_2294_n59272# A1 a_2030_n59272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2527 a_1634_n99458# a_1584_n66# a_1370_n99458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2528 GND A1 word24 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2529 a_2162_n43794# a_2112_n66# a_2030_n43794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2530 word642 A0 a_2162_n91364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2531 word893 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2532 GND A8 word201 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2533 GND A8 word762 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2534 a_446_n94914# A8 a_50_n94914# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2535 word519 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2536 word578 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2537 a_1898_n128284# a_1848_n66# a_1766_n128284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2538 a_2294_n141632# A1 a_1898_n141632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2539 a_2030_n12980# A2 a_1634_n12980# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2540 GND A7 word62 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2541 word571 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2542 GND A7 word887 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2543 VDD A7 a_528_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X2544 GND A7 word828 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2545 a_710_n86110# A7 a_446_n86110# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2546 word580 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2547 GND A9 word297 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2548 GND A3 word998 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2549 a_2030_n128568# A2 a_1634_n128568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2550 a_2294_n50184# A1 a_2030_n50184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2551 a_1634_n90370# a_1584_n66# a_1370_n90370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2552 GND A9 word238 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2553 a_2162_n144330# a_2112_n66# a_1898_n144330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2554 a_710_n16388# A7 a_446_n16388# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2555 GND A6 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2556 word106 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2557 a_2162_n59130# a_2112_n66# a_1898_n59130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2558 a_1634_n140070# a_1584_n66# a_1370_n140070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2559 GND A3 word896 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2560 word478 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2561 GND A1 word892 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2562 word29 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2563 a_710_n85684# A7 a_446_n85684# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2564 word559 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2565 word290 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2566 a_1370_n75602# a_1320_n66# a_1238_n75602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2567 word200 A0 a_2294_n28600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2568 a_2162_n67082# a_2112_n66# a_1898_n67082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2569 word620 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2570 a_974_n7442# A6 a_710_n7442# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2571 GND A5 word862 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2572 GND A6 word809 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2573 a_1106_n34422# a_1056_n66# a_842_n34422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2574 word683 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2575 word688 A0 a_2294_n97896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2576 GND A9 word504 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2577 a_710_n121610# A7 a_314_n121610# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2578 a_710_n54160# A7 a_314_n54160# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2579 GND A8 word25 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2580 a_2030_n27890# A2 a_1766_n27890# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2581 GND A5 word409 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2582 word495 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2583 word313 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2584 GND A5 word350 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2585 a_1238_n66088# A5 a_842_n66088# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2586 word676 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2587 a_2162_n112380# a_2112_n66# a_1898_n112380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2588 word243 a_2376_n66# a_2162_n34706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2589 GND A7 word98 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2590 a_2162_n27180# a_2112_n66# a_1898_n27180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2591 GND A9 word402 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2592 a_446_n31440# A8 a_182_n31440# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2593 a_2294_n65094# A1 a_2030_n65094# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2594 GND A8 word674 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2595 GND A9 word13 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2596 a_1370_n43652# a_1320_n66# a_1106_n43652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2597 GND A0 word996 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2598 word875 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2599 GND A8 word242 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2600 a_2162_n96476# a_2112_n66# a_1898_n96476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2601 word732 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2602 GND A7 word586 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2603 GND A8 word744 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2604 a_1766_n91222# A3 a_1502_n91222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2605 a_2294_n116640# A1 a_1898_n116640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2606 a_1766_n82844# A3 a_1502_n82844# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2607 GND A7 word44 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2608 a_1238_n122320# A5 a_842_n122320# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2609 GND A7 word869 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2610 word805 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2611 a_1370_n139644# a_1320_n66# a_1238_n139644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2612 a_2030_n74040# A2 a_1634_n74040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2613 a_1502_n101446# A4 a_1238_n101446# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2614 a_2030_n134390# A2 a_1766_n134390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2615 a_578_n136236# a_528_n66# a_314_n136236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2616 a_578_n127858# a_528_n66# a_314_n127858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2617 a_446_n6732# A8 a_182_n6732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2618 word28 A0 a_2294_n4176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2619 word62 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2620 a_446_n86252# A8 a_50_n86252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2621 a_1370_n12128# a_1320_n66# a_1238_n12128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2622 a_446_n77874# A8 a_50_n77874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2623 a_1766_n59982# A3 a_1502_n59982# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2624 GND A5 word967 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2625 word930 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2626 a_2294_n124592# A1 a_1898_n124592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2627 GND A0 word774 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2628 GND A7 word305 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2629 word77 a_2376_n66# a_2294_n11134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2630 word88 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2631 GND A1 word992 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2632 a_2294_n94488# A1 a_2030_n94488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2633 word861 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2634 GND A1 word933 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2635 a_1238_n130272# A5 a_974_n130272# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2636 a_1238_n121894# A5 a_842_n121894# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2637 a_2162_n2756# a_2112_n66# a_2030_n2756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2638 word937 a_2376_n66# a_2294_n133254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2639 a_1370_n81424# a_1320_n66# a_1106_n81424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2640 a_1370_n108120# a_1320_n66# a_1106_n108120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2641 a_2162_n127290# a_2112_n66# a_1898_n127290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2642 word939 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2643 a_1370_n130556# a_1320_n66# a_1238_n130556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2644 a_1766_n28458# A3 a_1502_n28458# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2645 GND A1 word501 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2646 GND A7 word361 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2647 a_974_n4886# A6 a_710_n4886# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2648 a_1766_n50894# A3 a_1502_n50894# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2649 GND A9 word59 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2650 a_1370_n58562# a_1320_n66# a_1238_n58562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2651 GND A7 word632 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2652 a_578_n104286# a_528_n66# a_446_n104286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2653 a_1370_n107694# a_1320_n66# a_1106_n107694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2654 a_1370_n116072# a_1320_n66# a_1106_n116072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2655 a_578_n23914# a_528_n66# a_446_n23914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2656 GND A5 word450 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2657 a_1106_n87104# a_1056_n66# a_842_n87104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2658 word910 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2659 a_1238_n137230# A5 a_842_n137230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2660 GND A2 word408 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2661 a_1106_n78726# a_1056_n66# a_974_n78726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2662 GND A6 word531 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2663 GND A4 word839 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2664 GND A7 word80 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2665 a_1106_n17382# a_1056_n66# a_842_n17382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2666 GND A1 word220 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2667 word684 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2668 GND A4 word997 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2669 a_1370_n27038# a_1320_n66# a_1106_n27038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2670 GND A0 word820 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2671 a_1766_n66230# A3 a_1370_n66230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2672 GND A7 word568 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2673 word966 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2674 word123 a_2376_n66# a_2162_n17666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2675 word714 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2676 word907 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2677 GND A3 word983 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2678 word831 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2679 a_446_n14400# A8 a_182_n14400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2680 word983 a_2376_n66# a_2162_n139786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2681 GND A8 word613 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2682 GND A8 word554 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2683 a_1370_n145466# a_1320_n66# a_1106_n145466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2684 word947 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2685 word611 a_2376_n66# a_2162_n86962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2686 GND A0 word876 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2687 GND A4 word775 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2688 a_578_n142058# a_528_n66# a_314_n142058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2689 a_578_n133680# a_528_n66# a_314_n133680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2690 a_50_n135952# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2691 a_446_n92074# A8 a_50_n92074# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2692 a_446_n83696# A8 a_50_n83696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2693 GND A6 word306 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2694 GND A3 word919 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2695 a_842_n118912# a_792_n66# a_710_n118912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2696 word919 a_2376_n66# a_2162_n130698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2697 a_710_n2472# A7 a_446_n2472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2698 a_50_n91932# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2699 word459 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2700 word725 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2701 a_842_n70916# a_792_n66# a_578_n70916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2702 word389 a_2376_n66# a_2294_n55438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2703 a_50_n104428# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2704 a_710_n119480# A7 a_314_n119480# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2705 a_1766_n34280# A3 a_1370_n34280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2706 GND A0 word308 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2707 GND A1 word325 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2708 GND A4 word301 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2709 GND A4 a_1320_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X2710 a_1898_n20222# a_1848_n66# a_1634_n20222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2711 GND A0 word206 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2712 a_182_n37404# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2713 a_1502_n19512# A4 a_1238_n19512# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2714 GND A6 word572 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2715 GND A5 word783 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2716 a_1898_n58704# a_1848_n66# a_1634_n58704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2717 a_1502_n113800# A4 a_1106_n113800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2718 a_710_n9430# A7 a_446_n9430# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2719 a_1766_n89092# A3 a_1370_n89092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2720 GND A3 word53 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2721 GND A4 word79 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2722 word655 a_2376_n66# a_2162_n93210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2723 a_842_n16530# a_792_n66# a_710_n16530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2724 GND A0 word574 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2725 word1007 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2726 GND A6 word411 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2727 word872 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2728 GND A1 word100 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2729 GND A0 word142 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2730 word813 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2731 word830 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2732 a_182_n1762# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2733 GND A4 word41 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2734 a_1502_n10424# A4 a_1238_n10424# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2735 a_842_n85826# a_792_n66# a_710_n85826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2736 a_1370_n93778# a_1320_n66# a_1238_n93778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2737 GND A8 word654 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2738 word988 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2739 GND A8 word595 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2740 a_50_n119338# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2741 GND A4 word76 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2742 GND A0 word472 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2743 word562 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2744 word794 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2745 a_50_n141774# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2746 word503 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2747 word798 A0 a_2162_n113516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2748 word31 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2749 GND A1 word588 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2750 word279 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2751 GND A6 word189 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2752 GND A5 word990 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2753 word496 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2754 GND A6 word130 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2755 word132 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2756 word191 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2757 a_1898_n35132# a_1848_n66# a_1766_n35132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2758 a_1106_n52598# a_1056_n66# a_842_n52598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2759 word401 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2760 a_842_n124734# a_792_n66# a_710_n124734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2761 a_50_n75318# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2762 word342 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2763 a_974_n92216# A6 a_578_n92216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2764 a_1106_n99458# a_1056_n66# a_974_n99458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2765 GND A2 word753 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2766 GND A6 word677 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2767 a_1502_n137088# A4 a_1238_n137088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2768 a_182_n8720# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2769 a_50_n110250# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2770 a_974_n22494# A6 a_578_n22494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2771 a_314_n64810# a_264_n66# a_182_n64810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2772 word396 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2773 a_50_n74892# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2774 a_842_n53876# a_792_n66# a_710_n53876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2775 word269 a_2376_n66# a_2294_n38398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2776 word4 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2777 word120 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2778 a_182_n43226# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2779 GND A0 word188 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2780 GND A4 word672 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2781 a_1106_n108404# a_1056_n66# a_842_n108404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2782 a_182_n34848# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2783 a_314_n72762# a_264_n66# a_182_n72762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2784 GND A8 word700 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2785 a_1106_n90370# a_1056_n66# a_842_n90370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2786 word398 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2787 word958 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2788 word899 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2789 a_1898_n64526# a_1848_n66# a_1766_n64526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2790 a_578_n21074# a_528_n66# a_446_n21074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2791 GND A3 word512 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2792 a_842_n101162# a_792_n66# a_578_n101162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2793 word176 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2794 GND A2 word960 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2795 a_974_n60266# A6 a_578_n60266# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2796 word610 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2797 word829 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2798 a_1370_n8862# a_1320_n66# a_1106_n8862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2799 a_578_n59556# a_528_n66# a_314_n59556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2800 a_842_n139644# a_792_n66# a_578_n139644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2801 a_314_n41238# a_264_n66# a_182_n41238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2802 a_974_n98748# A6 a_578_n98748# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2803 word662 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2804 VDD A1 a_2112_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X2805 word535 a_2376_n66# a_2162_n76170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2806 a_50_n125160# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2807 a_1634_n27322# a_1584_n66# a_1370_n27322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2808 GND A0 word454 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2809 GND A2 word1016 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2810 a_1766_n1194# A3 a_1502_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2811 a_182_n72620# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2812 a_1502_n54728# A4 a_1238_n54728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2813 word780 A0 a_2294_n110960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2814 word666 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2815 word379 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2816 word320 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2817 a_182_n11276# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2818 a_842_n68786# a_792_n66# a_578_n68786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2819 word173 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2820 word232 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2821 a_842_n108120# a_792_n66# a_578_n108120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2822 a_1898_n93920# a_1848_n66# a_1766_n93920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2823 a_1898_n32576# a_1848_n66# a_1766_n32576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2824 a_182_n49758# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2825 a_182_n58136# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2826 a_50_n81140# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2827 GND A3 word129 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2828 word383 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2829 a_314_n142342# a_264_n66# a_50_n142342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2830 word72 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2831 a_578_n97328# a_528_n66# a_446_n97328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2832 a_314_n133964# a_264_n66# a_50_n133964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2833 a_1898_n79436# a_1848_n66# a_1634_n79436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2834 GND A6 word659 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2835 word376 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2836 a_1238_n9572# A5 a_842_n9572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2837 a_1898_n18092# a_1848_n66# a_1634_n18092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2838 word153 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2839 GND A4 word225 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2840 a_842_n107694# a_792_n66# a_578_n107694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2841 word28 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2842 word437 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2843 a_974_n75176# A6 a_710_n75176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2844 word343 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2845 a_974_n134816# A6 a_578_n134816# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2846 a_1634_n56716# a_1584_n66# a_1502_n56716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2847 GND A4 word555 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2848 GND A6 word557 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2849 GND A0 word288 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2850 word959 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2851 a_314_n47770# a_264_n66# a_182_n47770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2852 a_314_n56148# a_264_n66# a_182_n56148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2853 word124 A0 a_2294_n17808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2854 a_1634_n106416# a_1584_n66# a_1502_n106416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2855 a_1106_n114226# a_1056_n66# a_974_n114226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2856 a_182_n40670# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2857 GND A2 word18 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2858 a_1106_n105848# a_1056_n66# a_842_n105848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2859 word439 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2860 GND A4 word69 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2861 word999 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2862 word112 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2863 word276 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2864 a_1898_n70348# a_1848_n66# a_1634_n70348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2865 a_1502_n78016# A4 a_1106_n78016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2866 word944 A0 a_2294_n134248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2867 word852 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2868 a_1502_n69638# A4 a_1106_n69638# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2869 GND A4 word552 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2870 a_182_n26186# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2871 word929 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2872 a_314_n110392# a_264_n66# a_50_n110392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2873 word870 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2874 word838 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2875 a_578_n57000# a_528_n66# a_314_n57000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2876 a_578_n65378# a_528_n66# a_314_n65378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2877 a_1898_n47486# a_1848_n66# a_1634_n47486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2878 a_842_n145466# a_792_n66# a_578_n145466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2879 a_50_n96050# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2880 a_1238_n46918# A5 a_842_n46918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2881 GND A3 word451 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2882 a_2294_n54302# A1 a_1898_n54302# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2883 word644 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2884 a_974_n111244# A6 a_710_n111244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2885 word768 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2886 GND A2 word840 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2887 a_1766_n114652# A3 a_1502_n114652# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2888 a_1634_n33144# a_1584_n66# a_1502_n33144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2889 word118 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2890 word317 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2891 word549 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2892 a_710_n42942# A7 a_314_n42942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2893 a_1634_n24766# a_1584_n66# a_1502_n24766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2894 GND A4 word330 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2895 a_1502_n60550# A4 a_1106_n60550# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2896 word926 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2897 a_1106_n143620# a_1056_n66# a_842_n143620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2898 a_1634_n135810# a_1584_n66# a_1370_n135810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2899 word23 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2900 GND A4 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2901 word542 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2902 word214 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2903 a_710_n89802# A7 a_446_n89802# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2904 a_2162_n15962# a_2112_n66# a_1898_n15962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2905 a_182_n55580# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2906 a_1502_n46066# A4 a_1238_n46066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2907 word446 A0 a_2162_n63532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2908 GND A7 word793 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2909 a_1502_n37688# A4 a_1238_n37688# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2910 a_314_n117350# a_264_n66# a_50_n117350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2911 word382 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2912 a_1898_n85258# a_1848_n66# a_1766_n85258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2913 a_710_n11418# A7 a_446_n11418# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2914 a_1898_n76880# a_1848_n66# a_1634_n76880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2915 word704 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2916 word957 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2917 GND A3 word658 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2918 word695 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2919 GND A3 word226 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2920 word975 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2921 GND A9 word101 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2922 a_2294_n22352# A1 a_1898_n22352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2923 a_710_n80714# A7 a_446_n80714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2924 a_2030_n62822# A2 a_1634_n62822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2925 a_2294_n13974# A1 a_2030_n13974# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2926 word224 A0 a_2294_n32008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2927 GND A5 word596 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2928 word1000 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2929 word998 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2930 a_710_n10992# A7 a_446_n10992# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2931 a_1238_n92642# A5 a_974_n92642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2932 a_1634_n103860# a_1584_n66# a_1370_n103860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2933 a_974_n117776# A6 a_710_n117776# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2934 GND A0 word600 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2935 GND A6 word774 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2936 a_1898_n138224# a_1848_n66# a_1634_n138224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2937 a_2030_n22920# A2 a_1766_n22920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2938 a_578_n71200# a_528_n66# a_314_n71200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2939 GND A3 word275 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2940 a_2294_n29310# A1 a_1898_n29310# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2941 GND A9 word367 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2942 a_2162_n22210# a_2112_n66# a_2030_n22210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2943 GND A3 word433 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2944 word487 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2945 GND A9 word308 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2946 word218 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2947 word809 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2948 a_710_n17950# A7 a_446_n17950# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2949 word299 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2950 word750 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2951 a_2030_n30872# A2 a_1634_n30872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2952 a_1238_n38256# A5 a_974_n38256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2953 word421 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2954 a_1238_n29878# A5 a_842_n29878# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2955 word489 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2956 a_2162_n91506# a_2112_n66# a_2030_n91506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2957 a_2294_n98606# A1 a_1898_n98606# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2958 GND A9 word206 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2959 word629 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2960 a_2162_n30162# a_2112_n66# a_2030_n30162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2961 a_2294_n37262# A1 a_1898_n37262# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2962 word360 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2963 a_2030_n77732# A2 a_1766_n77732# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2964 word197 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2965 word270 A0 a_2162_n38540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2966 word956 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2967 a_1634_n127148# a_1584_n66# a_1370_n127148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2968 a_1106_n126580# a_1056_n66# a_842_n126580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2969 word428 A0 a_2294_n60976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2970 a_2162_n68644# a_2112_n66# a_2030_n68644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2971 a_446_n72904# A8 a_50_n72904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2972 word423 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2973 GND A5 word149 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2974 GND A6 word820 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2975 GND A5 word90 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2976 a_1238_n20790# A5 a_974_n20790# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2977 word357 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2978 a_578_n108404# a_528_n66# a_446_n108404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2979 word694 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2980 a_2030_n37830# A2 a_1634_n37830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2981 word326 A0 a_2162_n46492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2982 GND A5 word479 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2983 GND A9 word142 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2984 GND A9 word83 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2985 word565 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2986 a_1238_n67650# A5 a_842_n67650# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2987 a_1238_n76028# A5 a_974_n76028# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2988 word687 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2989 word734 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2990 GND A9 word472 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2991 GND A9 word413 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2992 a_2294_n66656# A1 a_1898_n66656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2993 GND A3 word741 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2994 GND A1 word796 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2995 word323 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X2996 GND A1 word737 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2997 word741 a_2376_n66# a_2294_n105422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X2998 GND A9 word24 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X2999 a_1634_n45498# a_1584_n66# a_1370_n45498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3000 a_2030_n45782# A2 a_1766_n45782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3001 GND A5 word476 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3002 word878 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3003 a_1898_n144046# a_1848_n66# a_1766_n144046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3004 a_1370_n102724# a_1320_n66# a_1238_n102724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3005 a_446_n18518# A8 a_182_n18518# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3006 word592 A0 a_2294_n84264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3007 word690 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3008 word1001 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3009 a_2030_n14258# A2 a_1766_n14258# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3010 a_446_n87814# A8 a_50_n87814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3011 word158 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3012 word217 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3013 GND A5 word195 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3014 GND A7 word837 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3015 a_710_n79010# A7 a_446_n79010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3016 word931 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3017 GND A9 word247 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3018 a_1238_n140212# A5 a_842_n140212# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3019 GND A3 word948 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3020 a_1238_n131834# A5 a_974_n131834# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3021 a_1106_n8436# a_1056_n66# a_974_n8436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3022 GND A9 word188 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3023 a_1634_n83270# a_1584_n66# a_1502_n83270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3024 a_2030_n83554# A2 a_1634_n83554# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3025 GND A4 word801 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3026 a_1370_n21642# a_1320_n66# a_1238_n21642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3027 word997 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3028 GND A8 word87 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3029 a_2162_n74466# a_2112_n66# a_2030_n74466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3030 a_2294_n103008# A1 a_1898_n103008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3031 GND A1 word901 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3032 a_446_n105564# A8 a_50_n105564# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3033 GND A1 word512 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3034 a_1898_n112096# a_1848_n66# a_1766_n112096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3035 word240 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3036 a_710_n78584# A7 a_446_n78584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3037 GND A6 word16 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3038 a_1238_n100310# A5 a_842_n100310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3039 word983 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3040 a_1106_n41806# a_1056_n66# a_974_n41806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3041 a_1370_n126012# a_1320_n66# a_1106_n126012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3042 a_1370_n117634# a_1320_n66# a_1106_n117634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3043 GND A2 word89 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3044 a_578_n105848# a_528_n66# a_446_n105848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3045 GND A5 word520 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3046 word424 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3047 a_2294_n102582# A1 a_2030_n102582# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3048 a_710_n114510# A7 a_314_n114510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3049 GND A9 word454 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3050 a_1106_n27322# a_1056_n66# a_974_n27322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3051 a_2294_n72478# A1 a_1898_n72478# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3052 GND A8 word34 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3053 a_710_n47060# A7 a_314_n47060# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3054 GND A3 word723 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3055 word445 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3056 word626 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3057 word723 a_2376_n66# a_2162_n102866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3058 word193 a_2376_n66# a_2294_n27606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3059 word977 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3060 GND A1 word129 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3061 GND A4 word906 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3062 a_446_n24340# A8 a_182_n24340# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3063 a_710_n122462# A7 a_314_n122462# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3064 word1017 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3065 GND A8 word624 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3066 GND A2 word355 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3067 word681 a_2376_n66# a_2294_n96902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3068 GND A7 word536 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3069 GND A8 word753 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3070 GND A0 word946 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3071 word825 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3072 a_578_n143620# a_528_n66# a_314_n143620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3073 GND A8 word192 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3074 a_446_n93636# A8 a_50_n93636# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3075 a_1766_n75744# A3 a_1370_n75744# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3076 GND A1 word617 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3077 a_2294_n131976# A1 a_2030_n131976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3078 a_842_n9288# a_792_n66# a_710_n9288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3079 a_446_n32292# A8 a_182_n32292# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3080 GND A2 word194 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3081 GND A7 word819 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3082 GND A9 word288 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3083 a_578_n129136# a_528_n66# a_314_n129136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3084 a_1106_n5880# a_1056_n66# a_974_n5880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3085 word989 a_2376_n66# a_2294_n140638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3086 a_446_n79152# A8 a_50_n79152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3087 a_2030_n80998# A2 a_1634_n80998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3088 GND A0 word724 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3089 a_2162_n4034# a_2112_n66# a_2030_n4034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3090 a_974_n26612# A6 a_578_n26612# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3091 a_1766_n44220# A3 a_1370_n44220# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3092 word811 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3093 GND A3 word887 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3094 word887 a_2376_n66# a_2162_n126154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3095 word851 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3096 word526 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3097 word889 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3098 word792 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3099 a_1898_n4602# a_1848_n66# a_1634_n4602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3100 GND A7 word311 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3101 a_974_n6164# A6 a_710_n6164# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3102 a_50_n113942# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3103 a_1766_n43794# A3 a_1370_n43794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3104 GND A1 word392 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3105 GND A5 word853 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3106 GND A9 word495 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3107 a_1502_n132118# A4 a_1106_n132118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3108 a_1502_n123740# A4 a_1106_n123740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3109 GND A5 word794 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3110 a_1106_n24766# a_1056_n66# a_974_n24766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3111 a_1106_n33144# a_1056_n66# a_842_n33144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3112 GND A6 word151 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3113 a_1502_n109256# A4 a_1238_n109256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3114 word1018 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3115 GND A0 word212 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3116 GND A4 word1006 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3117 a_1766_n12270# A3 a_1370_n12270# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3118 GND A8 word665 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3119 GND A0 word770 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3120 GND A7 word577 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3121 GND A0 word928 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3122 a_1766_n5312# A3 a_1502_n5312# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3123 a_842_n34422# a_792_n66# a_578_n34422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3124 GND A8 word233 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3125 GND A7 word518 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3126 GND A8 word735 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3127 a_1238_n138082# A5 a_842_n138082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3128 word82 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3129 a_1370_n89234# a_1320_n66# a_1106_n89234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3130 GND A7 word35 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3131 a_446_n768# A8 a_182_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3132 GND A2 word235 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3133 a_1106_n62538# a_1056_n66# a_974_n62538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3134 a_1502_n100168# A4 a_1238_n100168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3135 GND A0 word826 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3136 word762 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3137 word412 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3138 word561 a_2376_n66# a_2294_n79862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3139 a_1370_n129988# a_1320_n66# a_1238_n129988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3140 a_446_n5454# A8 a_182_n5454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3141 a_50_n128852# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3142 GND A1 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3143 a_446_n76596# A8 a_50_n76596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3144 a_1766_n67082# A3 a_1370_n67082# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3145 GND A1 word556 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3146 word570 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3147 GND A5 word899 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3148 a_1502_n138650# A4 a_1238_n138650# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3149 GND A6 word256 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3150 word852 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3151 GND A3 word869 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3152 word409 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3153 a_1370_n80146# a_1320_n66# a_1106_n80146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3154 word869 a_2376_n66# a_2294_n123598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3155 a_50_n84832# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3156 word350 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3157 a_842_n63816# a_792_n66# a_578_n63816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3158 a_1370_n71768# a_1320_n66# a_1106_n71768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3159 a_1634_n6022# a_1584_n66# a_1502_n6022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3160 word339 a_2376_n66# a_2162_n48338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3161 GND A0 word258 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3162 word497 a_2376_n66# a_2294_n70774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3163 GND A7 word352 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3164 a_1370_n120900# a_1320_n66# a_1238_n120900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3165 GND A1 word492 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3166 GND A9 word50 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3167 a_1370_n57284# a_1320_n66# a_1238_n57284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3168 GND A1 word433 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3169 a_842_n49332# a_792_n66# a_710_n49332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3170 a_1238_n4602# A5 a_974_n4602# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3171 a_578_n31014# a_528_n66# a_446_n31014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3172 GND A7 word623 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3173 word822 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3174 a_578_n22636# a_528_n66# a_446_n22636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3175 word246 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3176 a_842_n102724# a_792_n66# a_578_n102724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3177 a_1766_n96476# A3 a_1502_n96476# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3178 GND A5 word30 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3179 word187 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3180 a_974_n61828# A6 a_578_n61828# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3181 a_1106_n77448# a_1056_n66# a_974_n77448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3182 GND A5 word733 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3183 GND A6 word522 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3184 a_1502_n115078# A4 a_1106_n115078# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3185 a_1502_n106700# A4 a_1106_n106700# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3186 a_578_n91932# a_528_n66# a_446_n91932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3187 word605 a_2376_n66# a_2294_n86110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3188 GND A0 word524 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3189 a_842_n31866# a_792_n66# a_578_n31866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3190 a_974_n38966# A6 a_710_n38966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3191 word957 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3192 a_1766_n2756# A3 a_1370_n2756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3193 GND A0 word92 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3194 word763 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3195 a_182_n21216# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3196 a_842_n87104# a_792_n66# a_710_n87104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3197 GND A4 word517 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3198 a_1370_n95056# a_1320_n66# a_1238_n95056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3199 a_182_n12838# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3200 a_314_n50752# a_264_n66# a_182_n50752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3201 a_50_n99742# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3202 word243 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3203 GND A8 word545 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3204 a_578_n60408# a_528_n66# a_314_n60408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3205 word661 a_2376_n66# a_2294_n94062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3206 a_1370_n144188# a_1320_n66# a_1106_n144188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3207 word803 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3208 a_842_n17382# a_792_n66# a_710_n17382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3209 a_50_n143052# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3210 word748 A0 a_2294_n106416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3211 a_446_n2898# A8 a_182_n2898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3212 a_50_n134674# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3213 a_314_n143904# a_264_n66# a_50_n143904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3214 word446 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3215 a_1898_n28032# a_1848_n66# a_1766_n28032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3216 a_1106_n45498# a_1056_n66# a_974_n45498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3217 GND A6 word297 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3218 a_842_n126012# a_792_n66# a_710_n126012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3219 a_710_n1194# A7 a_446_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3220 a_50_n90654# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3221 a_974_n76738# A6 a_710_n76738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3222 GND A5 word838 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3223 GND A0 word358 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3224 a_50_n103150# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3225 a_2294_n4886# A1 a_2030_n4886# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3226 a_182_n50610# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3227 a_314_n57710# a_264_n66# a_182_n57710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3228 GND A4 word134 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3229 a_1502_n32718# A4 a_1106_n32718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3230 GND A4 word292 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3231 word1010 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3232 a_842_n46776# a_792_n66# a_710_n46776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3233 word660 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3234 word863 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3235 GND A0 word138 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3236 GND A4 word622 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3237 a_182_n9572# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3238 a_182_n27748# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3239 a_182_n36126# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3240 a_314_n65662# a_264_n66# a_182_n65662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3241 a_314_n120332# a_264_n66# a_50_n120332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3242 word186 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3243 a_314_n111954# a_264_n66# a_50_n111954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3244 GND A6 word563 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3245 a_578_n66940# a_528_n66# a_314_n66940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3246 GND A4 word70 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3247 word54 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3248 word126 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3249 a_974_n112806# A6 a_710_n112806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3250 word223 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3251 a_974_n44788# A6 a_710_n44788# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3252 GND A6 word402 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3253 word560 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3254 word996 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3255 word804 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3256 word612 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3257 word745 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3258 word485 a_2376_n66# a_2294_n69070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3259 a_842_n84548# a_792_n66# a_710_n84548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3260 a_50_n118060# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3261 a_1502_n56006# A4 a_1238_n56006# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3262 GND A0 word404 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3263 GND A2 word907 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3264 a_182_n65520# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3265 a_50_n140496# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3266 a_1502_n47628# A4 a_1238_n47628# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3267 word435 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3268 word730 A0 a_2162_n103860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3269 word616 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3270 word22 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3271 GND A4 word397 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3272 word270 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3273 word182 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3274 word774 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3275 word428 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3276 word715 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3277 a_578_n34990# a_528_n66# a_446_n34990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3278 a_50_n74040# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3279 a_842_n123456# a_792_n66# a_710_n123456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3280 a_314_n135242# a_264_n66# a_50_n135242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3281 a_1106_n98180# a_1056_n66# a_974_n98180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3282 GND A6 word668 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3283 a_314_n126864# a_264_n66# a_50_n126864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3284 word326 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3285 a_1634_n11134# a_1584_n66# a_1502_n11134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3286 word103 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3287 word0 A0 a_2294_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3288 a_1502_n6874# A4 a_1106_n6874# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3289 GND A4 word175 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3290 a_1766_n139502# A3 a_1370_n139502# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3291 a_974_n127716# A6 a_578_n127716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3292 a_974_n59698# A6 a_578_n59698# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3293 GND A0 word670 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3294 a_842_n52598# a_792_n66# a_710_n52598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3295 a_1634_n49616# a_1584_n66# a_1370_n49616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3296 a_314_n49048# a_264_n66# a_182_n49048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3297 a_182_n33570# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3298 GND A2 word27 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3299 a_1502_n15678# A4 a_1106_n15678# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3300 a_1502_n24056# A4 a_1106_n24056# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3301 a_1106_n107126# a_1056_n66# a_842_n107126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3302 a_314_n71484# a_264_n66# a_182_n71484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3303 a_1370_n8010# a_1320_n66# a_1106_n8010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3304 word389 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3305 a_1634_n121752# a_1584_n66# a_1370_n121752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3306 word227 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3307 a_1898_n63248# a_1848_n66# a_1634_n63248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3308 word890 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3309 word540 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3310 GND A3 word562 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3311 word599 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3312 word894 A0 a_2162_n127148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3313 a_974_n200# A6 a_710_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3314 GND A3 word503 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3315 a_182_n19086# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3316 GND A0 word58 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3317 word68 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3318 a_1766_n130414# A3 a_1370_n130414# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3319 GND A3 word71 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3320 word229 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3321 word879 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3322 word820 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3323 a_578_n58278# a_528_n66# a_314_n58278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3324 a_1634_n40528# a_1584_n66# a_1370_n40528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3325 a_842_n138366# a_792_n66# a_578_n138366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3326 a_1370_n7584# a_1320_n66# a_1106_n7584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3327 a_1238_n39818# A5 a_974_n39818# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3328 word491 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3329 GND A3 word342 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3330 GND A3 word401 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3331 GND A4 word14 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3332 word127 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3333 a_2294_n38824# A1 a_2030_n38824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3334 a_842_n90370# a_792_n66# a_710_n90370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3335 a_974_n97470# A6 a_578_n97470# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3336 a_1766_n107552# A3 a_1370_n107552# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3337 a_2162_n31724# a_2112_n66# a_1898_n31724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3338 word267 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3339 a_1634_n17666# a_1584_n66# a_1370_n17666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3340 word876 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3341 word498 A0 a_2162_n70916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3342 word657 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3343 word655 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3344 a_1634_n128710# a_1584_n66# a_1502_n128710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3345 word741 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3346 a_1898_n107836# a_1848_n66# a_1766_n107836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3347 word434 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3348 word164 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3349 a_1238_n30730# A5 a_842_n30730# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3350 word427 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3351 a_842_n120900# a_792_n66# a_710_n120900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3352 a_182_n48480# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3353 word396 A0 a_2294_n56432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3354 GND A9 word212 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3355 a_314_n141064# a_264_n66# a_50_n141064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3356 GND A9 word153 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3357 a_1106_n144472# a_1056_n66# a_842_n144472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3358 a_578_n96050# a_528_n66# a_446_n96050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3359 a_314_n132686# a_264_n66# a_50_n132686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3360 a_1898_n78158# a_1848_n66# a_1766_n78158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3361 GND A6 word650 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3362 word652 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3363 GND A5 word216 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3364 GND A3 word608 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3365 GND A6 word946 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3366 GND A3 word176 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3367 word334 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3368 a_1766_n136946# A3 a_1502_n136946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3369 a_974_n133538# A6 a_578_n133538# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3370 a_710_n73614# A7 a_446_n73614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3371 word950 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3372 a_2162_n140212# a_2112_n66# a_2030_n140212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3373 a_2162_n131834# a_2112_n66# a_1898_n131834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3374 a_1238_n85542# A5 a_842_n85542# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3375 GND A4 word645 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3376 GND A2 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3377 a_2162_n46634# a_2112_n66# a_1898_n46634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3378 a_2162_n55012# a_2112_n66# a_2030_n55012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3379 word430 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3380 GND A0 word550 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3381 a_1502_n68360# A4 a_1106_n68360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3382 word662 A0 a_2162_n94204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3383 word539 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3384 word598 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3385 a_2162_n108972# a_2112_n66# a_1898_n108972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3386 GND A0 word40 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3387 GND A5 word324 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3388 word107 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3389 a_578_n64100# a_528_n66# a_314_n64100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3390 GND A5 word265 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3391 a_842_n144188# a_792_n66# a_578_n144188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3392 a_1238_n45640# A5 a_842_n45640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3393 GND A9 word317 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3394 GND A9 word258 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3395 a_2294_n44646# A1 a_2030_n44646# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3396 a_2294_n53024# A1 a_1898_n53024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3397 a_1634_n93210# a_1584_n66# a_1502_n93210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3398 word109 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3399 a_1766_n104996# A3 a_1502_n104996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3400 a_710_n41664# A7 a_314_n41664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3401 word249 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3402 a_710_n50042# A7 a_314_n50042# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3403 word14 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3404 GND A5 word321 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3405 GND A1 word912 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3406 word723 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3407 a_1238_n118912# A5 a_842_n118912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3408 a_1898_n113658# a_1848_n66# a_1634_n113658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3409 word310 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3410 a_710_n88524# A7 a_446_n88524# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3411 word597 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3412 a_2162_n14684# a_2112_n66# a_1898_n14684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3413 a_1634_n92784# a_1584_n66# a_1502_n92784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3414 GND A7 word784 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3415 word378 A0 a_2162_n53876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3416 word906 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3417 a_1634_n142484# a_1584_n66# a_1502_n142484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3418 word787 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3419 a_710_n10140# A7 a_446_n10140# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3420 word314 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3421 a_1766_n47912# A3 a_1370_n47912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3422 GND A6 word770 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3423 a_1238_n22068# A5 a_974_n22068# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3424 word307 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3425 word366 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3426 GND A6 word928 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3427 a_1238_n13690# A5 a_842_n13690# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3428 a_2030_n39108# A2 a_1766_n39108# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3429 word276 A0 a_2294_n39392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3430 word375 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3431 GND A9 word92 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3432 GND A1 word848 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3433 a_1634_n61260# a_1584_n66# a_1502_n61260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3434 word515 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3435 word793 a_2376_n66# a_2294_n112806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3436 a_2294_n12696# A1 a_2030_n12696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3437 a_2030_n61544# A2 a_1766_n61544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3438 GND A5 word587 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3439 a_2030_n121894# A2 a_1634_n121894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3440 a_2162_n115220# a_2112_n66# a_2030_n115220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3441 word696 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3442 word989 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3443 VDD A4 a_1320_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X3444 a_1238_n82986# A5 a_842_n82986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3445 a_1238_n91364# A5 a_974_n91364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3446 GND A6 word826 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3447 a_1766_n128284# A3 a_1502_n128284# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3448 a_2294_n81992# A1 a_2030_n81992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3449 a_974_n116498# A6 a_710_n116498# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3450 a_1634_n38398# a_1584_n66# a_1502_n38398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3451 word571 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3452 word644 A0 a_2294_n91648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3453 a_2162_n99316# a_2112_n66# a_2030_n99316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3454 word887 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3455 a_2162_n123172# a_2112_n66# a_2030_n123172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3456 a_1370_n104002# a_1320_n66# a_1238_n104002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3457 a_2162_n114794# a_2112_n66# a_1898_n114794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3458 a_2030_n30020# A2 a_1766_n30020# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3459 a_2162_n29594# a_2112_n66# a_1898_n29594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3460 word573 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3461 a_446_n33854# A8 a_182_n33854# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3462 word542 A0 a_2162_n77164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3463 GND A7 word889 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3464 GND A9 word358 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3465 GND A9 word299 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3466 word951 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3467 word48 A0 a_2294_n7016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3468 word478 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3469 word419 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3470 a_2294_n127432# A1 a_2030_n127432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3471 GND A5 word204 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3472 word108 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3473 a_1238_n28600# A5 a_842_n28600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3474 a_2294_n97328# A1 a_1898_n97328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3475 GND A3 word695 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3476 GND A1 word953 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3477 GND A7 word61 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3478 a_2162_n81850# a_2112_n66# a_1898_n81850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3479 a_2294_n88950# A1 a_2030_n88950# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3480 a_2162_n90228# a_2112_n66# a_2030_n90228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3481 word480 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3482 word822 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3483 word881 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3484 GND A9 word197 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3485 GND A3 word898 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3486 a_2030_n76454# A2 a_1634_n76454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3487 word638 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3488 GND A9 word138 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3489 GND A4 word751 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3490 a_710_n85968# A7 a_446_n85968# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3491 word1006 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3492 word862 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3493 GND A7 word381 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3494 word947 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3495 a_446_n80004# A8 a_50_n80004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3496 a_1766_n62112# A3 a_1370_n62112# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3497 GND A7 word322 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3498 a_974_n7726# A6 a_710_n7726# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3499 a_2162_n58988# a_2112_n66# a_1898_n58988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3500 GND A5 word140 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3501 word190 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3502 a_446_n10282# A8 a_182_n10282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3503 a_2162_n138082# a_2112_n66# a_2030_n138082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3504 GND A2 word98 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3505 a_1106_n34706# a_1056_n66# a_842_n34706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3506 a_578_n107126# a_528_n66# a_446_n107126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3507 word956 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3508 word678 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3509 word315 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3510 word725 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3511 word66 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3512 GND A2 word586 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3513 GND A9 word404 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3514 a_1238_n101162# A5 a_842_n101162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3515 GND A1 word728 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3516 a_1502_n141632# A4 a_1106_n141632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3517 a_2294_n57000# A1 a_2030_n57000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3518 GND A9 word15 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3519 word395 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3520 a_1370_n43936# a_1320_n66# a_1106_n43936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3521 word869 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3522 GND A0 word998 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3523 GND A8 word244 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3524 a_1766_n91506# A3 a_1502_n91506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3525 word734 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3526 a_1238_n139644# A5 a_842_n139644# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3527 a_446_n17240# A8 a_182_n17240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3528 word301 a_2376_n66# a_2294_n42942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3529 a_710_n115362# A7 a_314_n115362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3530 a_1766_n30162# A3 a_1370_n30162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3531 GND A1 word237 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3532 GND A7 word97 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3533 GND A1 word296 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3534 word701 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3535 GND A0 word896 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3536 GND A2 word305 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3537 word631 a_2376_n66# a_2162_n89802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3538 a_1502_n101730# A4 a_1238_n101730# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3539 a_1502_n110108# A4 a_1238_n110108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3540 a_1370_n139928# a_1320_n66# a_1238_n139928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3541 a_578_n136520# a_528_n66# a_314_n136520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3542 word30 A0 a_2162_n4460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3543 word933 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3544 a_446_n86536# A8 a_50_n86536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3545 a_1766_n68644# A3 a_1502_n68644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3546 a_2294_n133254# A1 a_2030_n133254# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3547 a_446_n25192# A8 a_182_n25192# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3548 GND A1 word21 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3549 word90 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3550 GND A2 word203 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3551 GND A7 word769 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3552 word922 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3553 a_1106_n7158# a_1056_n66# a_974_n7158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3554 word79 a_2376_n66# a_2162_n11418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3555 word863 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3556 a_1238_n130556# A5 a_974_n130556# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3557 GND A2 word361 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3558 a_2030_n82276# A2 a_1766_n82276# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3559 word939 a_2376_n66# a_2162_n133538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3560 a_578_n144472# a_528_n66# a_314_n144472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3561 a_710_n5312# A7 a_446_n5312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3562 word479 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3563 a_1370_n81708# a_1320_n66# a_1106_n81708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3564 word61 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3565 word637 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3566 a_842_n12412# a_792_n66# a_710_n12412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3567 a_1370_n11986# a_1320_n66# a_1238_n11986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3568 a_974_n19512# A6 a_578_n19512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3569 word567 a_2376_n66# a_2162_n80714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3570 GND A2 word632 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3571 GND A2 word691 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3572 word988 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3573 a_1370_n130840# a_1320_n66# a_1238_n130840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3574 GND A3 word837 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3575 a_1766_n37120# A3 a_1502_n37120# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3576 GND A8 word78 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3577 GND A7 word363 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3578 a_2162_n73188# a_2112_n66# a_2030_n73188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3579 GND A1 word833 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3580 a_446_n104286# A8 a_50_n104286# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3581 word837 a_2376_n66# a_2294_n119054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3582 a_1370_n58846# a_1320_n66# a_1238_n58846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3583 a_1370_n67224# a_1320_n66# a_1238_n67224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3584 GND A6 word7 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3585 GND A2 word80 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3586 word476 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3587 a_1370_n107978# a_1320_n66# a_1106_n107978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3588 GND A8 word566 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3589 a_1370_n116356# a_1320_n66# a_1106_n116356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3590 GND A1 word401 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3591 GND A7 word261 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3592 a_578_n104570# a_528_n66# a_446_n104570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3593 a_50_n106842# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3594 a_1766_n36694# A3 a_1502_n36694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3595 GND A2 word410 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3596 a_1502_n125018# A4 a_1106_n125018# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3597 a_1106_n26044# a_1056_n66# a_974_n26044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3598 GND A9 word445 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3599 a_1106_n17666# a_1056_n66# a_842_n17666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3600 a_2294_n71200# A1 a_1898_n71200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3601 GND A2 word568 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3602 word254 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3603 word125 a_2376_n66# a_2294_n17950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3604 GND A0 word162 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3605 GND A2 word466 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3606 a_1106_n86962# a_1056_n66# a_842_n86962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3607 word968 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3608 a_182_n4602# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3609 GND A1 word120 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3610 a_2030_n97186# A2 a_1634_n97186# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3611 GND A4 word897 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3612 a_1502_n124592# A4 a_1106_n124592# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3613 a_710_n121184# A7 a_314_n121184# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3614 word1008 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3615 GND A8 word615 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3616 GND A4 word96 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3617 a_1370_n35274# a_1320_n66# a_1106_n35274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3618 word949 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3619 a_1370_n26896# a_1320_n66# a_1106_n26896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3620 GND A8 word183 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3621 GND A7 word527 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3622 GND A0 word878 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3623 a_50_n144614# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3624 a_446_n92358# A8 a_50_n92358# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3625 GND A1 word608 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3626 a_2162_n88098# a_2112_n66# a_2030_n88098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3627 a_2030_n2614# A2 a_1766_n2614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3628 word91 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3629 a_446_n83980# A8 a_50_n83980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3630 GND A1 word176 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3631 GND A2 word185 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3632 GND A6 word308 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3633 GND A8 word671 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3634 a_710_n2756# A7 a_446_n2756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3635 word520 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3636 GND A5 word908 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3637 word86 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3638 a_974_n25334# A6 a_578_n25334# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3639 GND A2 word673 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3640 GND A2 word931 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3641 word802 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3642 GND A3 word819 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3643 word581 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3644 word819 a_2376_n66# a_2162_n116498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3645 GND A4 word362 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3646 a_50_n77732# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3647 a_1898_n20506# a_1848_n66# a_1634_n20506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3648 a_1370_n122178# a_1320_n66# a_1238_n122178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3649 a_50_n121042# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3650 a_1898_n3324# a_1848_n66# a_1766_n3324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3651 GND A0 word208 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3652 word447 a_2376_n66# a_2162_n63674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3653 GND A7 word302 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3654 a_50_n112664# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3655 GND A5 word844 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3656 GND A4 word201 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3657 GND A6 word574 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3658 word291 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3659 GND A5 word785 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3660 word831 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3661 a_1106_n23488# a_1056_n66# a_974_n23488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3662 GND A6 word142 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3663 a_1766_n89376# A3 a_1370_n89376# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3664 a_842_n104002# a_792_n66# a_578_n104002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3665 word772 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3666 a_1502_n1904# A4 a_1238_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3667 a_446_n98890# A8 a_50_n98890# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3668 a_974_n63106# A6 a_578_n63106# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3669 word225 a_2376_n66# a_2294_n32150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3670 word293 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3671 a_974_n54728# A6 a_578_n54728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3672 GND A6 word413 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3673 GND A2 word507 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3674 word1009 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3675 word874 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3676 GND A0 word144 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3677 GND A2 word706 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3678 GND A4 word938 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3679 word815 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3680 GND A4 word43 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3681 a_1502_n10708# A4 a_1238_n10708# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3682 word555 a_2376_n66# a_2162_n79010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3683 word990 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3684 word855 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3685 a_1766_n342# A3 a_1502_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3686 a_842_n33144# a_792_n66# a_578_n33144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3687 word191 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3688 GND A0 word474 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3689 GND A2 word977 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3690 word37 a_2376_n66# a_2294_n5454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3691 word132 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3692 word505 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3693 GND A1 word649 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3694 word708 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3695 word686 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3696 GND A7 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3697 a_1766_n80288# A3 a_1370_n80288# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3698 a_182_n14116# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3699 word498 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3700 word871 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3701 a_314_n43652# a_264_n66# a_182_n43652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3702 a_1106_n61260# a_1056_n66# a_974_n61260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3703 word193 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3704 word888 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3705 a_1370_n2614# a_1320_n66# a_1238_n2614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3706 a_446_n4176# A8 a_182_n4176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3707 a_50_n127574# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3708 a_1898_n9856# a_1848_n66# a_1766_n9856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3709 word403 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3710 GND A1 word488 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3711 word856 A0 a_2294_n121752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3712 a_314_n136804# a_264_n66# a_50_n136804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3713 GND A2 word755 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3714 GND A6 word679 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3715 word681 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3716 word396 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3717 a_974_n22778# A6 a_578_n22778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3718 GND A6 word188 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3719 a_974_n78016# A6 a_710_n78016# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3720 a_50_n83554# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3721 word398 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3722 a_182_n43510# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3723 a_578_n99742# a_528_n66# a_446_n99742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3724 GND A4 word674 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3725 GND A2 word752 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3726 GND A2 word811 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3727 a_1238_n3324# A5 a_974_n3324# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3728 a_842_n48054# a_792_n66# a_710_n48054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3729 a_1898_n64810# a_1848_n66# a_1766_n64810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3730 GND A7 word614 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3731 a_842_n101446# a_792_n66# a_578_n101446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3732 word813 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3733 a_182_n29026# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3734 a_578_n21358# a_528_n66# a_446_n21358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3735 word178 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3736 a_314_n58562# a_264_n66# a_182_n58562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3737 a_182_n51462# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3738 GND A3 word82 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3739 a_974_n60550# A6 a_578_n60550# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3740 a_314_n113232# a_264_n66# a_50_n113232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3741 GND A6 word513 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3742 a_578_n59840# a_528_n66# a_314_n59840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3743 a_578_n68218# a_528_n66# a_314_n68218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3744 word456 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3745 a_842_n139928# a_792_n66# a_578_n139928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3746 word63 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3747 a_1898_n72762# a_1848_n66# a_1634_n72762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3748 word666 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3749 word173 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3750 a_974_n37688# A6 a_710_n37688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3751 GND A2 word1018 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3752 word19 a_2376_n66# a_2162_n2898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3753 a_842_n30588# a_792_n66# a_578_n30588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3754 word946 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3755 word43 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3756 a_578_n67792# a_528_n66# a_314_n67792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3757 word754 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3758 a_182_n11560# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3759 a_50_n98464# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3760 GND A4 word449 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3761 a_1370_n85400# a_1320_n66# a_1238_n85400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3762 a_2162_n18802# a_2112_n66# a_2030_n18802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3763 word234 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3764 a_1634_n96902# a_1584_n66# a_1502_n96902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3765 word735 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3766 a_182_n58420# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3767 a_50_n133396# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3768 a_1898_n32860# a_1848_n66# a_1766_n32860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3769 word444 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3770 word343 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3771 a_314_n142626# a_264_n66# a_50_n142626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3772 word724 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3773 word437 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3774 word74 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3775 word378 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3776 a_578_n36268# a_528_n66# a_446_n36268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3777 a_1238_n9856# A5 a_842_n9856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3778 GND A6 word288 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3779 a_578_n27890# a_528_n66# a_446_n27890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3780 GND A5 word286 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3781 a_842_n107978# a_792_n66# a_578_n107978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3782 a_182_n66372# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3783 word30 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3784 GND A3 word246 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3785 a_182_n57994# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3786 a_50_n80998# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3787 a_2294_n16814# A1 a_1898_n16814# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3788 word439 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3789 a_974_n75460# A6 a_710_n75460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3790 a_314_n119764# a_264_n66# a_50_n119764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3791 a_314_n128142# a_264_n66# a_50_n128142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3792 GND A6 word559 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3793 word276 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3794 a_1634_n2188# a_1584_n66# a_1502_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3795 word1020 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3796 a_710_n13832# A7 a_446_n13832# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3797 GND A0 word290 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3798 word721 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3799 a_1106_n114510# a_1056_n66# a_974_n114510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3800 GND A0 word620 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3801 word278 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3802 word854 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3803 a_182_n8294# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3804 word219 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3805 a_1634_n64952# a_1584_n66# a_1502_n64952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3806 GND A4 word554 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3807 GND A4 word613 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3808 a_182_n26470# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3809 a_314_n64384# a_264_n66# a_182_n64384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3810 a_314_n110676# a_264_n66# a_50_n110676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3811 word118 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3812 a_1898_n47770# a_1848_n66# a_1634_n47770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3813 word497 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3814 word45 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3815 GND A0 word676 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3816 GND A3 word35 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3817 word111 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3818 GND A3 word453 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3819 a_1502_n77874# A4 a_1106_n77874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3820 word1002 A0 a_2162_n142484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3821 GND A6 word791 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3822 a_1766_n123314# A3 a_1502_n123314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3823 a_4876_164# A7 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X3824 a_974_n111528# A6 a_710_n111528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3825 word483 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3826 word214 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3827 a_1634_n33428# a_1584_n66# a_1502_n33428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3828 a_710_n51604# A7 a_314_n51604# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3829 word770 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3830 GND A5 word391 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3831 word928 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3832 word987 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3833 a_842_n83270# a_792_n66# a_710_n83270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3834 GND A4 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3835 a_2162_n33002# a_2112_n66# a_1898_n33002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3836 a_1502_n46350# A4 a_1238_n46350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3837 word826 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3838 word13 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3839 word443 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3840 word448 A0 a_2294_n63816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3841 a_1898_n109114# a_1848_n66# a_1634_n109114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3842 word607 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3843 GND A4 word388 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3844 word959 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3845 word377 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3846 word436 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3847 GND A3 word660 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3848 word900 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3849 a_842_n122178# a_792_n66# a_710_n122178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3850 word346 A0 a_2162_n49332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3851 GND A9 word162 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3852 a_182_n72194# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3853 GND A3 word228 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3854 GND A9 word103 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3855 a_2030_n140212# A2 a_1634_n140212# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3856 a_2294_n31014# A1 a_2030_n31014# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3857 a_314_n125586# a_264_n66# a_50_n125586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3858 word661 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3859 a_1634_n129562# a_1584_n66# a_1502_n129562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3860 a_1238_n92926# A5 a_974_n92926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3861 GND A6 word896 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3862 a_1502_n5596# A4 a_1106_n5596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3863 a_1238_n31582# A5 a_842_n31582# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3864 a_1898_n100026# a_1848_n66# a_1634_n100026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3865 a_1766_n129846# A3 a_1370_n129846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3866 word319 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3867 word501 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3868 a_1634_n39960# a_1584_n66# a_1370_n39960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3869 word641 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3870 GND A4 word654 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3871 a_1898_n138508# a_1848_n66# a_1634_n138508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3872 a_1502_n14400# A4 a_1106_n14400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3873 word282 A0 a_2162_n40244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3874 a_2030_n100310# A2 a_1766_n100310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3875 word751 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3876 word218 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3877 a_1634_n120474# a_1584_n66# a_1502_n120474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3878 word159 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3879 a_1766_n25902# A3 a_1370_n25902# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3880 word612 A0 a_2294_n87104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3881 word421 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3882 GND A3 word435 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3883 a_1502_n83696# A4 a_1238_n83696# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3884 a_1502_n92074# A4 a_1238_n92074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3885 word220 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3886 a_2294_n60408# A1 a_2030_n60408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3887 a_1766_n120758# A3 a_1370_n120758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3888 GND A5 word274 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3889 word482 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3890 a_842_n137088# a_792_n66# a_578_n137088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3891 a_1238_n38540# A5 a_974_n38540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3892 GND A9 word267 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3893 a_1634_n86110# a_1584_n66# a_1370_n86110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3894 GND A9 word208 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3895 word199 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3896 word1017 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3897 GND A5 word271 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3898 word357 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3899 a_2162_n77306# a_2112_n66# a_1898_n77306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3900 a_2162_n101162# a_2112_n66# a_1898_n101162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3901 word732 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3902 a_1238_n46492# A5 a_842_n46492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3903 a_446_n108404# A8 a_50_n108404# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3904 a_1898_n106558# a_1848_n66# a_1634_n106558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3905 word606 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3906 GND A5 word210 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3907 a_446_n20222# A8 a_182_n20222# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3908 GND A6 word36 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3909 a_1634_n85684# a_1584_n66# a_1370_n85684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3910 word687 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3911 a_2162_n139644# a_2112_n66# a_1898_n139644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3912 a_446_n11844# A8 a_182_n11844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3913 a_2030_n115220# A2 a_1634_n115220# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3914 GND A2 word64 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3915 word328 A0 a_2294_n46776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3916 word485 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3917 GND A9 word144 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3918 a_1106_n143194# a_1056_n66# a_842_n143194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3919 word323 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3920 word737 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3921 a_1634_n135384# a_1584_n66# a_1370_n135384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3922 a_2294_n105422# A1 a_1898_n105422# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3923 word316 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3924 GND A3 word599 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3925 GND A6 word937 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3926 GND A9 word474 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3927 a_2294_n75318# A1 a_2030_n75318# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3928 a_1238_n111102# A5 a_974_n111102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3929 a_1766_n144046# A3 a_1370_n144046# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3930 word325 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3931 a_1238_n102724# A5 a_842_n102724# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3932 GND A3 word743 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3933 a_974_n132260# A6 a_578_n132260# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3934 a_1634_n54160# a_1584_n66# a_1370_n54160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3935 word465 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3936 word743 a_2376_n66# a_2162_n105706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3937 a_2030_n123172# A2 a_1766_n123172# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3938 GND A5 word537 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3939 word441 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3940 a_1238_n84264# A5 a_842_n84264# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3941 a_1898_n144330# a_1848_n66# a_1766_n144330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3942 a_2162_n130556# a_2112_n66# a_1898_n130556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3943 a_1238_n75886# A5 a_974_n75886# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3944 a_710_n125302# A7 a_314_n125302# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3945 a_2162_n36978# a_2112_n66# a_2030_n36978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3946 a_2162_n45356# a_2112_n66# a_1898_n45356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3947 a_710_n116924# A7 a_314_n116924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3948 a_974_n109398# A6 a_710_n109398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3949 a_710_n49474# A7 a_314_n49474# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3950 GND A8 word51 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3951 word521 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3952 word594 A0 a_2162_n84548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3953 word837 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3954 word1003 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3955 word530 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3956 a_2294_n134816# A1 a_1898_n134816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3957 a_446_n26754# A8 a_182_n26754# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3958 a_446_n35132# A8 a_182_n35132# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3959 GND A7 word839 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3960 GND A1 word32 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3961 GND A1 word1005 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3962 a_1106_n8720# a_1056_n66# a_974_n8720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3963 a_2030_n92216# A2 a_1634_n92216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3964 GND A9 word249 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3965 word901 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3966 a_2294_n43368# A1 a_2030_n43368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3967 a_1766_n112096# A3 a_1370_n112096# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3968 a_2294_n34990# A1 a_1898_n34990# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3969 word100 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3970 a_1370_n21926# a_1320_n66# a_1238_n21926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3971 a_710_n40386# A7 a_314_n40386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3972 a_1370_n30304# a_1320_n66# a_1238_n30304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3973 GND A8 word89 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3974 GND A8 word148 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3975 word831 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3976 word714 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3977 word216 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3978 a_446_n105848# A8 a_50_n105848# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3979 word772 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3980 a_2030_n138082# A2 a_1634_n138082# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3981 a_1898_n112380# a_1848_n66# a_1766_n112380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3982 a_710_n78868# A7 a_446_n78868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3983 a_710_n87246# A7 a_446_n87246# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3984 word588 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3985 GND A1 word141 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3986 a_2162_n145466# a_2112_n66# a_1898_n145466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3987 GND A6 word18 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3988 GND A7 word775 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3989 GND A8 word636 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3990 GND A7 word272 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3991 GND A7 word331 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3992 word897 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3993 a_1370_n117918# a_1320_n66# a_1106_n117918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3994 a_974_n9004# A6 a_710_n9004# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3995 a_1766_n55012# A3 a_1502_n55012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3996 GND A1 word412 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X3997 GND A8 word706 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X3998 a_1766_n46634# A3 a_1502_n46634# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X3999 word37 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4000 GND A3 word640 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4001 GND A7 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4002 GND A6 word919 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4003 GND A3 word784 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4004 a_1766_n141490# A3 a_1502_n141490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4005 word906 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4006 GND A1 word780 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4007 word265 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4008 GND A5 word578 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4009 word628 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4010 GND A5 word519 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4011 GND A2 word536 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4012 a_1106_n96902# a_1056_n66# a_974_n96902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4013 GND A4 word967 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4014 a_2162_n51178# a_2112_n66# a_1898_n51178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4015 a_2294_n58278# A1 a_2030_n58278# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4016 a_710_n122746# A7 a_314_n122746# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4017 word345 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4018 a_1370_n45214# a_1320_n66# a_1106_n45214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4019 GND A8 word33 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4020 GND A8 word253 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4021 GND A8 word755 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4022 GND A0 word948 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4023 GND A8 word194 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4024 a_2162_n89660# a_2112_n66# a_1898_n89660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4025 word251 a_2376_n66# a_2162_n35842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4026 a_446_n93920# A8 a_50_n93920# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4027 a_1766_n84406# A3 a_1370_n84406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4028 a_1898_n127290# a_1848_n66# a_1634_n127290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4029 GND A7 word55 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4030 GND A7 word106 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4031 a_2294_n140638# A1 a_1898_n140638# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4032 a_446_n32576# A8 a_182_n32576# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4033 a_1766_n14684# A3 a_1502_n14684# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4034 a_1766_n23062# A3 a_1502_n23062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4035 word564 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4036 GND A7 word880 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4037 GND A9 word21 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4038 a_578_n129420# a_528_n66# a_314_n129420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4039 GND A9 word290 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4040 word883 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4041 a_446_n79436# A8 a_50_n79436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4042 GND A8 word752 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4043 a_2294_n117776# A1 a_1898_n117776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4044 a_446_n18092# A8 a_182_n18092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4045 GND A7 word52 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4046 word872 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4047 GND A1 word944 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4048 GND A1 word885 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4049 word813 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4050 word889 a_2376_n66# a_2294_n126438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4051 a_710_n84690# A7 a_446_n84690# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4052 a_2030_n75176# A2 a_1766_n75176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4053 a_578_n137372# a_528_n66# a_314_n137372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4054 a_578_n128994# a_528_n66# a_314_n128994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4055 GND A4 word742 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4056 word853 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4057 a_1370_n13264# a_1320_n66# a_1238_n13264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4058 word587 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4059 word938 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4060 word794 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4061 GND A0 word782 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4062 GND A7 word313 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4063 GND A7 word372 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4064 word517 a_2376_n66# a_2294_n73614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4065 a_50_n122604# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4066 GND A1 word453 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4067 a_974_n6448# A6 a_710_n6448# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4068 a_1766_n52456# A3 a_1370_n52456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4069 GND A5 word855 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4070 word19 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4071 a_2162_n3892# a_2112_n66# a_2030_n3892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4072 a_1106_n33428# a_1056_n66# a_842_n33428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4073 GND A6 word153 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4074 word1006 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4075 GND A8 word516 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4076 a_1370_n131692# a_1320_n66# a_1238_n131692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4077 word365 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4078 a_1502_n109540# A4 a_1238_n109540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4079 GND A9 word395 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4080 GND A2 word577 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4081 a_1502_n131976# A4 a_1106_n131976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4082 word204 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4083 a_842_n34706# a_792_n66# a_578_n34706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4084 GND A8 word235 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4085 GND A7 word579 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4086 a_1238_n138366# A5 a_842_n138366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4087 GND A0 word112 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4088 word351 a_2376_n66# a_2162_n50042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4089 GND A2 word416 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4090 a_1106_n79862# a_1056_n66# a_974_n79862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4091 GND A1 word660 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4092 a_1238_n129988# A5 a_974_n129988# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4093 GND A7 word88 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4094 a_1370_n89518# a_1320_n66# a_1106_n89518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4095 a_710_n114084# A7 a_314_n114084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4096 word941 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4097 GND A1 word228 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4098 word958 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4099 a_50_n137514# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4100 GND A8 word133 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4101 GND A0 word828 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4102 a_446_n5738# A8 a_182_n5738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4103 word55 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4104 a_446_n85258# A8 a_50_n85258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4105 a_446_n76880# A8 a_50_n76880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4106 GND A7 word576 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4107 GND A5 word960 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4108 a_2294_n123598# A1 a_1898_n123598# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4109 word140 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4110 GND A6 word317 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4111 GND A8 word621 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4112 GND A1 word985 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4113 GND A3 word930 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4114 GND A2 word352 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4115 GND A6 word258 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4116 a_1106_n70774# a_1056_n66# a_842_n70774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4117 word854 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4118 a_1238_n120900# A5 a_842_n120900# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4119 a_710_n4034# A7 a_446_n4034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4120 a_578_n62822# a_528_n66# a_314_n62822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4121 a_1370_n80430# a_1320_n66# a_1106_n80430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4122 GND A4 word783 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4123 a_578_n143194# a_528_n66# a_314_n143194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4124 a_2294_n7726# A1 a_1898_n7726# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4125 word52 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4126 word569 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4127 GND A2 word682 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4128 a_842_n11134# a_792_n66# a_710_n11134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4129 a_1634_n6306# a_1584_n66# a_1502_n6306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4130 GND A7 word354 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4131 GND A2 word881 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4132 word531 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4133 GND A3 word769 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4134 word769 a_2376_n66# a_2294_n109398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4135 a_842_n49616# a_792_n66# a_710_n49616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4136 a_1370_n57568# a_1320_n66# a_1238_n57568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4137 GND A7 word625 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4138 word830 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4139 word733 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4140 a_578_n22920# a_528_n66# a_446_n22920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4141 a_1898_n13406# a_1848_n66# a_1634_n13406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4142 word397 a_2376_n66# a_2294_n56574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4143 word988 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4144 a_50_n105564# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4145 word248 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4146 a_182_n61402# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4147 a_314_n68502# a_264_n66# a_182_n68502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4148 GND A1 word333 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4149 GND A6 word524 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4150 GND A5 word735 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4151 a_1106_n16388# a_1056_n66# a_842_n16388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4152 a_1898_n82702# a_1848_n66# a_1766_n82702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4153 a_578_n30872# a_528_n66# a_446_n30872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4154 a_974_n56006# A6 a_578_n56006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4155 word175 a_2376_n66# a_2162_n25050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4156 word959 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4157 GND A0 word94 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4158 GND A2 word457 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4159 word900 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4160 word824 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4161 word765 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4162 a_182_n3324# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4163 a_1370_n95340# a_1320_n66# a_1238_n95340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4164 word663 a_2376_n66# a_2162_n94346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4165 a_842_n17666# a_792_n66# a_710_n17666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4166 a_50_n143336# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4167 word717 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4168 a_50_n134958# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4169 a_2030_n1336# A2 a_1634_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4170 a_1766_n73188# A3 a_1502_n73188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4171 a_446_n91080# A8 a_50_n91080# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4172 GND A1 word540 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4173 GND A0 word582 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4174 GND A4 word417 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4175 a_1502_n72904# A4 a_1238_n72904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4176 a_314_n36552# a_264_n66# a_182_n36552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4177 word448 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4178 word821 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4179 a_1106_n54160# a_1056_n66# a_842_n54160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4180 a_1898_n28316# a_1848_n66# a_1766_n28316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4181 GND A6 word299 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4182 a_842_n86962# a_792_n66# a_710_n86962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4183 a_1898_n50752# a_1848_n66# a_1766_n50752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4184 a_710_n1478# A7 a_446_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4185 a_182_n67934# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4186 a_50_n90938# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4187 a_314_n129704# a_264_n66# a_50_n129704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4188 word511 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4189 GND A5 word840 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4190 word806 A0 a_2162_n114652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4191 word346 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4192 a_1634_n3750# a_1584_n66# a_1370_n3750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4193 word77 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4194 a_974_n24056# A6 a_578_n24056# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4195 GND A0 word360 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4196 GND A2 word664 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4197 a_1898_n97612# a_1848_n66# a_1634_n97612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4198 GND A2 word922 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4199 a_1502_n9714# A4 a_1238_n9714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4200 GND A6 word138 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4201 word572 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4202 word791 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4203 GND A4 word353 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4204 a_50_n76454# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4205 GND A4 word294 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4206 word348 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4207 a_1370_n63390# a_1320_n66# a_1106_n63390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4208 a_974_n93352# A6 a_578_n93352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4209 word924 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4210 a_1898_n2046# a_1848_n66# a_1634_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4211 GND A2 word761 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4212 a_182_n9856# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4213 a_182_n36410# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4214 a_50_n111386# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4215 a_1502_n18518# A4 a_1238_n18518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4216 a_314_n65946# a_264_n66# a_182_n65946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4217 GND A4 word192 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4218 a_1106_n132402# a_1056_n66# a_974_n132402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4219 a_314_n120616# a_264_n66# a_50_n120616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4220 GND A6 word565 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4221 word282 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4222 word910 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4223 a_1898_n57710# a_1848_n66# a_1766_n57710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4224 word560 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4225 word181 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4226 a_1502_n87814# A4 a_1106_n87814# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4227 a_182_n44362# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4228 a_1106_n69070# a_1056_n66# a_842_n69070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4229 a_182_n35984# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4230 word284 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4231 GND A6 word404 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4232 word1000 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4233 word998 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4234 word406 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4235 word966 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4236 word865 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4237 a_1898_n65662# a_1848_n66# a_1634_n65662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4238 word907 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4239 GND A4 word34 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4240 word182 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4241 word645 a_2376_n66# a_2294_n91790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4242 word896 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4243 GND A2 word968 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4244 a_50_n140780# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4245 a_1634_n42942# a_1584_n66# a_1502_n42942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4246 GND A1 word640 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4247 word618 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4248 word677 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4249 GND A4 word399 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4250 GND A4 word458 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4251 a_314_n42374# a_264_n66# a_182_n42374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4252 word86 A0 a_2162_n12412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4253 word184 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4254 a_974_n99884# A6 a_578_n99884# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4255 a_1898_n25760# a_1848_n66# a_1766_n25760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4256 a_1898_n34138# a_1848_n66# a_1634_n34138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4257 a_842_n123740# a_792_n66# a_710_n123740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4258 a_50_n126296# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4259 a_1502_n55864# A4 a_1238_n55864# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4260 a_1502_n64242# A4 a_1238_n64242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4261 a_314_n135526# a_264_n66# a_50_n135526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4262 GND A6 word670 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4263 word672 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4264 word387 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4265 word328 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4266 a_1634_n11418# a_1584_n66# a_1502_n11418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4267 a_974_n21500# A6 a_578_n21500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4268 a_578_n29168# a_528_n66# a_446_n29168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4269 a_2030_n11702# A2 a_1766_n11702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4270 GND A3 word196 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4271 a_182_n59272# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4272 a_50_n82276# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4273 word389 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4274 a_50_n73898# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4275 GND A0 word240 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4276 a_578_n98464# a_528_n66# a_446_n98464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4277 GND A2 word802 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4278 a_1502_n24340# A4 a_1106_n24340# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4279 a_1106_n107410# a_1056_n66# a_842_n107410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4280 a_314_n71768# a_264_n66# a_182_n71768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4281 a_1634_n10992# a_1584_n66# a_1502_n10992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4282 GND A4 word233 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4283 a_1238_n2046# A5 a_974_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4284 a_974_n135952# A6 a_578_n135952# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4285 word804 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4286 a_578_n20080# a_528_n66# a_446_n20080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4287 a_1766_n9288# A3 a_1502_n9288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4288 word491 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4289 a_842_n100168# a_792_n66# a_578_n100168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4290 a_182_n19370# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4291 a_182_n50184# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4292 a_314_n57284# a_264_n66# a_182_n57284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4293 GND A0 word60 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4294 word132 A0 a_2294_n18944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4295 a_1502_n32292# A4 a_1106_n32292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4296 a_1106_n115362# a_1056_n66# a_974_n115362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4297 GND A2 word26 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4298 word127 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4299 GND A6 word445 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4300 a_1106_n106984# a_1056_n66# a_842_n106984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4301 word506 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4302 a_842_n138650# a_792_n66# a_578_n138650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4303 a_1370_n7868# a_1320_n66# a_1106_n7868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4304 GND A0 word626 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4305 word447 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4306 word1007 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4307 GND A3 word403 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4308 a_1898_n71484# a_1848_n66# a_1766_n71484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4309 a_1502_n79152# A4 a_1106_n79152# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4310 word655 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4311 word657 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4312 word952 A0 a_2294_n135384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4313 a_1766_n116214# A3 a_1370_n116214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4314 a_1766_n107836# A3 a_1370_n107836# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4315 a_710_n44504# A7 a_314_n44504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4316 word164 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4317 a_1634_n26328# a_1584_n66# a_1370_n26328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4318 a_2030_n26612# A2 a_1634_n26612# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4319 word937 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4320 GND A2 word1009 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4321 word34 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4322 a_1634_n17950# a_1584_n66# a_1370_n17950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4323 GND A5 word341 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4324 word427 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4325 word878 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4326 word659 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4327 word743 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4328 a_1238_n56432# A5 a_974_n56432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4329 a_2162_n102724# a_2112_n66# a_2030_n102724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4330 a_50_n97186# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4331 word225 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4332 word617 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4333 a_2162_n17524# a_2112_n66# a_2030_n17524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4334 word652 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4335 word398 A0 a_2162_n56716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4336 word557 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4337 a_1502_n70064# A4 a_1106_n70064# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4338 a_314_n141348# a_264_n66# a_50_n141348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4339 a_1634_n145324# a_1584_n66# a_1370_n145324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4340 a_1106_n144756# a_1056_n66# a_842_n144756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4341 word334 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4342 a_314_n132970# a_264_n66# a_50_n132970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4343 word369 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4344 word909 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4345 a_1898_n17098# a_1848_n66# a_1766_n17098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4346 GND A3 word610 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4347 a_842_n106700# a_792_n66# a_578_n106700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4348 GND A6 word948 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4349 GND A9 word112 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4350 a_182_n65094# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4351 GND A3 word178 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4352 word430 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4353 GND A7 word801 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4354 a_2030_n133112# A2 a_1634_n133112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4355 a_2294_n15536# A1 a_1898_n15536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4356 a_314_n118486# a_264_n66# a_50_n118486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4357 GND A6 word550 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4358 a_1898_n86394# a_1848_n66# a_1634_n86394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4359 a_1238_n94204# A5 a_974_n94204# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4360 a_710_n12554# A7 a_446_n12554# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4361 a_1238_n85826# A5 a_842_n85826# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4362 a_2294_n84832# A1 a_1898_n84832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4363 word451 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4364 word105 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4365 word269 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4366 a_1634_n72052# a_1584_n66# a_1370_n72052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4367 word591 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4368 word983 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4369 word845 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4370 a_1634_n63674# a_1584_n66# a_1370_n63674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4371 a_2162_n126012# a_2112_n66# a_1898_n126012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4372 a_2162_n117634# a_2112_n66# a_2030_n117634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4373 word232 A0 a_2294_n33144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4374 GND A4 word545 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4375 a_1634_n113374# a_1584_n66# a_1370_n113374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4376 a_1766_n18802# A3 a_1502_n18802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4377 word161 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4378 GND A6 word782 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4379 word102 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4380 GND A3 word385 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4381 a_974_n110250# A6 a_710_n110250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4382 a_2030_n32434# A2 a_1766_n32434# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4383 a_710_n50326# A7 a_314_n50326# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4384 a_710_n41948# A7 a_314_n41948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4385 word919 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4386 word286 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4387 a_1898_n122320# a_1848_n66# a_1634_n122320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4388 word535 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4389 a_1634_n79010# a_1584_n66# a_1502_n79010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4390 a_2162_n23346# a_2112_n66# a_2030_n23346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4391 a_710_n88808# A7 a_446_n88808# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4392 word226 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4393 word307 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4394 word967 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4395 a_1238_n39392# A5 a_974_n39392# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4396 a_1634_n142768# a_1584_n66# a_1502_n142768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4397 word375 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4398 a_2162_n92642# a_2112_n66# a_2030_n92642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4399 a_2294_n99742# A1 a_1898_n99742# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4400 a_1898_n130272# a_1848_n66# a_1766_n130272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4401 a_2294_n112806# A1 a_2030_n112806# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4402 a_446_n13122# A8 a_182_n13122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4403 word950 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4404 word368 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4405 a_1634_n78584# a_1584_n66# a_1502_n78584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4406 GND A7 word17 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4407 word278 A0 a_2162_n39676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4408 a_2030_n108120# A2 a_1634_n108120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4409 GND A9 word94 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4410 a_1106_n136094# a_1056_n66# a_974_n136094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4411 a_578_n132402# a_528_n66# a_314_n132402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4412 a_2294_n21358# A1 a_1898_n21358# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4413 a_2030_n61828# A2 a_1766_n61828# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4414 GND A5 word648 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4415 word698 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4416 word85 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4417 GND A5 word589 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4418 GND A3 word549 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4419 a_1238_n91648# A5 a_974_n91648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4420 GND A6 word828 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4421 GND A5 word157 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4422 a_2294_n59840# A1 a_1898_n59840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4423 a_1238_n104002# A5 a_842_n104002# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4424 GND A1 word748 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4425 a_2162_n52740# a_2112_n66# a_2030_n52740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4426 word415 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4427 a_2294_n90654# A1 a_1898_n90654# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4428 word492 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4429 word702 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4430 a_2030_n116072# A2 a_1766_n116072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4431 a_2030_n38966# A2 a_1766_n38966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4432 a_1634_n47060# a_1584_n66# a_1502_n47060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4433 word573 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4434 word889 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4435 a_1238_n77164# A5 a_974_n77164# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4436 word742 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4437 a_1898_n137230# a_1848_n66# a_1766_n137230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4438 word214 A0 a_2162_n30588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4439 GND A7 word117 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4440 a_710_n118202# A7 a_314_n118202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4441 GND A9 word421 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4442 word150 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4443 a_1766_n33002# A3 a_1502_n33002# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4444 a_710_n109824# A7 a_314_n109824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4445 word634 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4446 a_2162_n60692# a_2112_n66# a_2030_n60692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4447 word471 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4448 a_2294_n67792# A1 a_1898_n67792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4449 word575 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4450 word544 A0 a_2294_n77448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4451 GND A9 word360 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4452 GND A9 word32 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4453 word953 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4454 a_1898_n145182# a_1848_n66# a_1634_n145182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4455 word751 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4456 a_446_n28032# A8 a_182_n28032# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4457 a_578_n100452# a_528_n66# a_446_n100452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4458 word638 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4459 a_446_n19654# A8 a_182_n19654# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4460 GND A1 word41 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4461 GND A5 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4462 word110 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4463 GND A9 word199 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4464 GND A2 word322 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4465 GND A4 word812 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4466 a_578_n138934# a_528_n66# a_314_n138934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4467 a_2030_n76738# A2 a_1634_n76738# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4468 GND A9 word357 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4469 a_2030_n15394# A2 a_1634_n15394# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4470 GND A8 word98 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4471 word949 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4472 word1008 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4473 a_2162_n67650# a_2112_n66# a_2030_n67650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4474 a_446_n107126# A8 a_50_n107126# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4475 a_2162_n76028# a_2112_n66# a_1898_n76028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4476 a_1898_n105280# a_1848_n66# a_1766_n105280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4477 a_446_n10566# A8 a_182_n10566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4478 GND A6 word27 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4479 word762 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4480 a_578_n107410# a_528_n66# a_446_n107410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4481 GND A8 word586 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4482 a_2162_n129988# a_2112_n66# a_2030_n129988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4483 word1017 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4484 a_1766_n39534# A3 a_1370_n39534# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4485 a_2294_n104144# A1 a_1898_n104144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4486 word680 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4487 word17 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4488 word68 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4489 GND A9 word465 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4490 a_2294_n74040# A1 a_2030_n74040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4491 a_1238_n101446# A5 a_842_n101446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4492 a_1502_n141916# A4 a_1106_n141916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4493 a_1766_n134390# A3 a_1370_n134390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4494 GND A1 word789 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4495 a_1106_n42942# a_1056_n66# a_974_n42942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4496 GND A2 word97 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4497 a_2030_n44788# A2 a_1634_n44788# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4498 a_578_n106984# a_528_n66# a_446_n106984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4499 GND A5 word528 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4500 GND A5 word469 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4501 a_1106_n89802# a_1056_n66# a_842_n89802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4502 a_1238_n139928# A5 a_842_n139928# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4503 a_2162_n120900# a_2112_n66# a_2030_n120900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4504 a_1502_n127432# A4 a_1238_n127432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4505 a_710_n124024# A7 a_314_n124024# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4506 a_1766_n30446# A3 a_1370_n30446# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4507 a_2162_n35700# a_2112_n66# a_2030_n35700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4508 GND A8 word42 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4509 a_710_n115646# A7 a_314_n115646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4510 a_710_n48196# A7 a_314_n48196# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4511 a_1370_n29736# a_1320_n66# a_1238_n29736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4512 GND A8 word203 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4513 GND A0 word898 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4514 word271 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4515 word935 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4516 word201 a_2376_n66# a_2294_n28742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4517 a_446_n86820# A8 a_50_n86820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4518 a_1766_n68928# A3 a_1502_n68928# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4519 word792 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4520 GND A1 word196 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4521 a_446_n25476# A8 a_182_n25476# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4522 GND A1 word137 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4523 GND A7 word830 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4524 GND A8 word691 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4525 a_1106_n80714# a_1056_n66# a_974_n80714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4526 word924 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4527 GND A8 word632 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4528 GND A9 word240 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4529 a_1238_n130840# A5 a_974_n130840# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4530 GND A2 word363 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4531 GND A8 word761 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4532 word833 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4533 a_578_n144756# a_528_n66# a_314_n144756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4534 a_2294_n119054# A1 a_1898_n119054# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4535 a_446_n94772# A8 a_50_n94772# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4536 word639 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4537 a_1370_n20648# a_1320_n66# a_1238_n20648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4538 word990 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4539 GND A8 word80 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4540 GND A3 word839 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4541 GND A1 word505 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4542 a_446_n104570# A8 a_50_n104570# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4543 GND A3 word997 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4544 word839 a_2376_n66# a_2162_n119338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4545 GND A2 word202 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4546 a_710_n77590# A7 a_446_n77590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4547 a_2030_n59698# A2 a_1766_n59698# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4548 a_1370_n67508# a_1320_n66# a_1238_n67508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4549 word921 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4550 word997 a_2376_n66# a_2294_n141774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4551 GND A1 word73 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4552 GND A6 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4553 word537 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4554 a_2162_n144188# a_2112_n66# a_1898_n144188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4555 word467 a_2376_n66# a_2162_n66514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4556 GND A0 word732 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4557 GND A8 word568 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4558 a_1370_n116640# a_1320_n66# a_1106_n116640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4559 a_50_n115504# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4560 GND A7 word263 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4561 a_1766_n36978# A3 a_1502_n36978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4562 word690 A0 a_2162_n98180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4563 a_1106_n17950# a_1056_n66# a_842_n17950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4564 a_1106_n26328# a_1056_n66# a_974_n26328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4565 GND A6 word162 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4566 GND A3 word775 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4567 word775 a_2376_n66# a_2162_n110250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4568 word619 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4569 GND A1 word69 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4570 a_1106_n95624# a_1056_n66# a_974_n95624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4571 word970 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4572 GND A9 word345 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4573 GND A5 word861 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4574 a_1502_n133254# A4 a_1106_n133254# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4575 GND A4 word899 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4576 a_1502_n124876# A4 a_1106_n124876# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4577 a_710_n121468# A7 a_314_n121468# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4578 word1010 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4579 a_842_n27606# a_792_n66# a_578_n27606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4580 a_1370_n35558# a_1320_n66# a_1106_n35558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4581 GND A8 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4582 GND A7 word529 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4583 GND A8 word185 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4584 a_4876_164# A7 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X4585 word93 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4586 word891 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4587 a_446_n31298# A8 a_182_n31298# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4588 GND A8 word673 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4589 word931 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4590 a_446_n7016# A8 a_182_n7016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4591 a_446_n78158# A8 a_50_n78158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4592 GND A7 word526 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4593 GND A5 word910 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4594 a_974_n25618# A6 a_578_n25618# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4595 GND A6 word267 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4596 a_1106_n72052# a_1056_n66# a_842_n72052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4597 word804 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4598 GND A3 word880 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4599 a_1238_n122178# A5 a_842_n122178# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4600 a_578_n55722# a_528_n66# a_314_n55722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4601 a_1106_n63674# a_1056_n66# a_974_n63674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4602 a_578_n136094# a_528_n66# a_314_n136094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4603 word785 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4604 a_974_n94914# A6 a_578_n94914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4605 GND A0 word714 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4606 GND A5 word966 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4607 GND A5 word907 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4608 a_50_n121326# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4609 word449 a_2376_n66# a_2294_n63958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4610 GND A7 word304 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4611 a_974_n5170# A6 a_710_n5170# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4612 a_50_n112948# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4613 a_1766_n51178# A3 a_1502_n51178# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4614 GND A1 word385 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4615 GND A1 word444 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4616 GND A4 word262 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4617 a_1370_n81282# a_1320_n66# a_1106_n81282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4618 word293 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4619 a_1106_n32150# a_1056_n66# a_842_n32150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4620 a_842_n64952# a_792_n66# a_578_n64952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4621 a_1766_n98038# A3 a_1370_n98038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4622 GND A6 word144 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4623 word347 a_2376_n66# a_2162_n49474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4624 word146 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4625 a_1766_n89660# A3 a_1370_n89660# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4626 word706 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4627 word991 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4628 word938 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4629 a_182_n54302# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4630 GND A0 word266 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4631 a_182_n45924# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4632 a_1106_n79010# a_1056_n66# a_974_n79010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4633 GND A4 word999 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4634 GND A4 word940 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4635 a_578_n23772# a_528_n66# a_446_n23772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4636 a_842_n33428# a_792_n66# a_578_n33428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4637 GND A7 word570 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4638 a_1766_n626# A3 a_1502_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4639 word39 a_2376_n66# a_2162_n5738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4640 a_1106_n78584# a_1056_n66# a_974_n78584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4641 word909 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4642 a_1238_n137088# A5 a_842_n137088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4643 GND A7 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4644 word283 a_2376_n66# a_2162_n40386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4645 a_974_n62964# A6 a_578_n62964# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4646 GND A4 word838 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4647 a_314_n52314# a_264_n66# a_182_n52314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4648 word932 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4649 a_314_n43936# a_264_n66# a_182_n43936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4650 word683 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4651 word890 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4652 word613 a_2376_n66# a_2294_n87246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4653 word755 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4654 a_50_n136236# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4655 word405 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4656 GND A7 word350 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4657 GND A0 word532 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4658 GND A1 word549 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4659 a_446_n4460# A8 a_182_n4460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4660 a_50_n127858# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4661 a_1502_n65804# A4 a_1238_n65804# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4662 a_1766_n66088# A3 a_1370_n66088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4663 word398 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4664 a_182_n22352# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4665 a_182_n13974# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4666 word251 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4667 word845 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4668 a_578_n61544# a_528_n66# a_314_n61544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4669 a_842_n141632# a_792_n66# a_578_n141632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4670 word811 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4671 a_182_n69212# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4672 a_50_n92216# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4673 word756 A0 a_2294_n107552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4674 a_50_n83838# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4675 GND A3 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4676 a_2294_n6448# A1 a_1898_n6448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4677 GND A0 word310 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4678 GND A2 word872 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4679 word741 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4680 word522 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4681 GND A4 word303 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4682 word47 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4683 a_842_n48338# a_792_n66# a_710_n48338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4684 a_1238_n3608# A5 a_974_n3608# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4685 a_578_n30020# a_528_n66# a_446_n30020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4686 a_1898_n12128# a_1848_n66# a_1766_n12128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4687 a_842_n70774# a_792_n66# a_578_n70774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4688 a_974_n77874# A6 a_710_n77874# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4689 word815 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4690 a_842_n101730# a_792_n66# a_578_n101730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4691 a_182_n29310# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4692 a_182_n60124# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4693 a_314_n67224# a_264_n66# a_182_n67224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4694 a_50_n104286# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4695 word180 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4696 GND A0 word366 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4697 a_1106_n125302# a_1056_n66# a_842_n125302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4698 a_182_n51746# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4699 a_314_n58846# a_264_n66# a_182_n58846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4700 a_1502_n33854# A4 a_1106_n33854# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4701 a_1502_n42232# A4 a_1106_n42232# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4702 a_314_n113516# a_264_n66# a_50_n113516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4703 GND A6 word515 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4704 a_1106_n116924# a_1056_n66# a_974_n116924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4705 GND A0 word696 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4706 GND A3 word55 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4707 a_1898_n81424# a_1848_n66# a_1634_n81424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4708 word1018 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4709 GND A5 word81 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4710 word1022 A0 a_2162_n145324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4711 word871 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4712 a_182_n28884# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4713 a_182_n37262# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4714 word950 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4715 word948 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4716 a_182_n2046# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4717 GND A6 word571 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4718 a_710_n9288# A7 a_446_n9288# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4719 a_50_n98748# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4720 a_842_n86110# a_792_n66# a_710_n86110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4721 GND A3 word52 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4722 GND A4 word78 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4723 word74 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4724 word595 a_2376_n66# a_2162_n84690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4725 a_842_n16388# a_792_n66# a_710_n16388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4726 a_50_n133680# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4727 a_50_n142058# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4728 word627 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4729 a_974_n113942# A6 a_710_n113942# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4730 a_1634_n35842# a_1584_n66# a_1370_n35842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4731 a_314_n142910# a_264_n66# a_50_n142910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4732 word439 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4733 a_1502_n10282# A4 a_1238_n10282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4734 word134 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4735 a_1898_n27038# a_1848_n66# a_1634_n27038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4736 GND A6 word290 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4737 a_842_n85684# a_792_n66# a_710_n85684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4738 a_842_n125018# a_792_n66# a_710_n125018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4739 a_50_n119196# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4740 word344 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4741 word502 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4742 a_182_n66656# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4743 a_314_n128426# a_264_n66# a_50_n128426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4744 word738 A0 a_2162_n104996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4745 word337 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4746 word278 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4747 a_1898_n96334# a_1848_n66# a_1766_n96334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4748 word782 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4749 word563 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4750 word723 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4751 a_842_n124592# a_792_n66# a_710_n124592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4752 a_50_n75176# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4753 a_842_n54160# a_792_n66# a_710_n54160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4754 word462 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4755 a_974_n92074# A6 a_578_n92074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4756 GND A6 word676 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4757 GND A0 word190 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4758 GND A4 word615 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4759 a_182_n8578# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4760 word111 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4761 word1019 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4762 a_314_n64668# a_264_n66# a_182_n64668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4763 word179 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4764 a_1634_n114936# a_1584_n66# a_1502_n114936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4765 a_314_n110960# a_264_n66# a_50_n110960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4766 a_974_n128852# A6 a_578_n128852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4767 word231 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4768 GND A0 word678 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4769 word172 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4770 GND A3 word455 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4771 a_1502_n86536# A4 a_1106_n86536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4772 word1004 A0 a_2294_n142768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4773 GND A6 word793 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4774 word119 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4775 a_182_n43084# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4776 word667 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4777 a_1106_n108262# a_1056_n66# a_842_n108262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4778 a_2030_n102724# A2 a_1766_n102724# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4779 a_1370_n9146# a_1320_n66# a_1106_n9146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4780 GND A6 word395 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4781 word397 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4782 word989 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4783 a_1898_n64384# a_1848_n66# a_1766_n64384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4784 a_1238_n63816# A5 a_842_n63816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4785 word605 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4786 word607 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4787 word902 A0 a_2162_n128284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4788 a_2162_n24908# a_2112_n66# a_1898_n24908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4789 a_2294_n62822# A1 a_2030_n62822# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4790 GND A0 word66 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4791 a_710_n37404# A7 a_314_n37404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4792 a_2030_n19512# A2 a_1634_n19512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4793 a_1634_n50042# a_1584_n66# a_1370_n50042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4794 word237 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4795 word887 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4796 word828 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4797 word668 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4798 word377 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4799 a_2162_n104002# a_2112_n66# a_2030_n104002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4800 word609 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4801 word15 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4802 a_1238_n49332# A5 a_842_n49332# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4803 GND A4 word390 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4804 a_314_n41096# a_264_n66# a_182_n41096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4805 a_842_n69070# a_792_n66# a_578_n69070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4806 word175 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4807 word661 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4808 word1020 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4809 a_1898_n131834# a_1848_n66# a_1634_n131834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4810 a_1634_n88524# a_1584_n66# a_1502_n88524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4811 GND A3 word289 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4812 word348 A0 a_2294_n49616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4813 a_1634_n138224# a_1584_n66# a_1502_n138224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4814 a_182_n72478# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4815 GND A3 word230 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4816 a_314_n125870# a_264_n66# a_50_n125870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4817 a_314_n134248# a_264_n66# a_50_n134248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4818 word663 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4819 word12 A0 a_2294_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4820 word155 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4821 a_2294_n22920# A1 a_2030_n22920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4822 a_1898_n108972# a_1848_n66# a_1634_n108972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4823 word319 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4824 a_2030_n10424# A2 a_1634_n10424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4825 word442 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4826 GND A3 word560 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4827 a_1502_n5880# A4 a_1106_n5880# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4828 GND A6 word898 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4829 GND A3 word128 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4830 a_1238_n31866# A5 a_842_n31866# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4831 a_1238_n40244# A5 a_974_n40244# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4832 word380 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4833 word503 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4834 a_2030_n117634# A2 a_1634_n117634# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4835 word643 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4836 a_2294_n30872# A1 a_2030_n30872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4837 word71 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4838 a_578_n97186# a_528_n66# a_446_n97186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4839 a_1898_n79294# a_1848_n66# a_1634_n79294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4840 word211 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4841 word284 A0 a_2294_n40528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4842 a_314_n70490# a_264_n66# a_182_n70490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4843 a_2162_n39818# a_2112_n66# a_1898_n39818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4844 GND A9 word491 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4845 word342 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4846 a_974_n134674# A6 a_578_n134674# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4847 word541 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4848 a_1634_n56574# a_1584_n66# a_1502_n56574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4849 a_1502_n92358# A4 a_1238_n92358# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4850 word182 A0 a_2162_n26044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4851 a_1502_n83980# A4 a_1238_n83980# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4852 a_1634_n106274# a_1584_n66# a_1502_n106274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4853 a_1106_n114084# a_1056_n66# a_974_n114084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4854 word484 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4855 word438 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4856 a_1502_n69496# A4 a_1106_n69496# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4857 a_2162_n30730# a_2112_n66# a_1898_n30730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4858 word120 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4859 a_2294_n37830# A1 a_2030_n37830# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4860 a_2294_n46208# A1 a_1898_n46208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4861 GND A9 word427 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4862 a_710_n43226# A7 a_314_n43226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4863 a_1634_n25050# a_1584_n66# a_1502_n25050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4864 word547 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4865 word606 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4866 GND A2 word1000 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4867 a_2030_n25334# A2 a_1766_n25334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4868 GND A5 word332 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4869 word869 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4870 word236 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4871 GND A5 word273 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4872 word650 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4873 word734 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4874 a_1238_n46776# A5 a_842_n46776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4875 a_1238_n55154# A5 a_974_n55154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4876 word485 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4877 word608 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4878 GND A9 word266 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4879 a_446_n20506# A8 a_182_n20506# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4880 a_2294_n45782# A1 a_2030_n45782# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4881 a_1634_n85968# a_1584_n66# a_1370_n85968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4882 word257 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4883 a_314_n140070# a_264_n66# a_50_n140070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4884 a_1106_n143478# a_1056_n66# a_842_n143478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4885 a_1634_n135668# a_1584_n66# a_1370_n135668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4886 word645 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4887 a_1898_n114794# a_1848_n66# a_1766_n114794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4888 word318 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4889 GND A7 word851 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4890 GND A6 word939 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4891 a_1766_n144330# A3 a_1370_n144330# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4892 GND A7 word792 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4893 a_2030_n63106# A2 a_1634_n63106# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4894 a_2030_n54728# A2 a_1766_n54728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4895 GND A5 word539 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4896 GND A5 word598 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4897 a_710_n11276# A7 a_446_n11276# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4898 a_1238_n84548# A5 a_842_n84548# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4899 a_2162_n54018# a_2112_n66# a_2030_n54018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4900 GND A3 word657 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4901 a_974_n118060# A6 a_710_n118060# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4902 GND A8 word53 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4903 word383 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4904 GND A1 word856 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4905 GND A3 word801 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4906 a_710_n49758# A7 a_314_n49758# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4907 word523 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4908 word839 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4909 word801 a_2376_n66# a_2294_n113942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4910 a_710_n80572# A7 a_446_n80572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4911 a_2162_n107978# a_2112_n66# a_1898_n107978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4912 word1005 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4913 a_2162_n116356# a_2112_n66# a_2030_n116356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4914 word164 A0 a_2294_n23488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4915 word997 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4916 word862 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4917 a_446_n35416# A8 a_182_n35416# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4918 GND A9 word41 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4919 GND A9 word310 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4920 word903 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4921 a_2294_n52030# A1 a_1898_n52030# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4922 word652 A0 a_2294_n92784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4923 a_1766_n112380# A3 a_1370_n112380# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4924 word647 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4925 a_710_n40670# A7 a_314_n40670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4926 a_2030_n31156# A2 a_1634_n31156# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4927 GND A1 word905 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4928 GND A2 word331 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4929 a_2162_n22068# a_2112_n66# a_2030_n22068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4930 a_2294_n29168# A1 a_1898_n29168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4931 GND A2 word272 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4932 a_2030_n69638# A2 a_1634_n69638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4933 a_710_n87530# A7 a_446_n87530# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4934 a_1502_n105422# A4 a_1106_n105422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4935 word590 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4936 word991 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4937 GND A9 word366 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4938 GND A9 word307 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4939 a_2030_n129988# A2 a_1766_n129988# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4940 word56 A0 a_2294_n8152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4941 a_2162_n13690# a_2112_n66# a_1898_n13690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4942 a_1370_n16104# a_1320_n66# a_1106_n16104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4943 word958 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4944 word430 A0 a_2162_n61260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4945 word899 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4946 a_2294_n98464# A1 a_1898_n98464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4947 GND A8 word708 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4948 GND A1 word961 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4949 a_2162_n6732# a_2112_n66# a_1898_n6732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4950 a_2162_n82986# a_2112_n66# a_1898_n82986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4951 word488 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4952 a_2162_n91364# a_2112_n66# a_2030_n91364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4953 a_2294_n111528# A1 a_2030_n111528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4954 word39 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4955 word359 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4956 GND A7 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4957 word300 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4958 GND A8 word536 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4959 GND A9 word85 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4960 a_2294_n20080# A1 a_1898_n20080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4961 a_1370_n134532# a_1320_n66# a_1106_n134532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4962 a_2030_n120900# A2 a_1766_n120900# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4963 a_578_n131124# a_528_n66# a_314_n131124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4964 word689 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4965 a_2030_n60550# A2 a_1634_n60550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4966 GND A5 word580 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4967 word630 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4968 a_974_n8862# A6 a_710_n8862# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4969 GND A9 word415 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4970 GND A6 word819 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4971 GND A2 word106 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4972 a_1106_n35842# a_1056_n66# a_842_n35842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4973 a_2030_n46066# A2 a_1766_n46066# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4974 a_578_n108262# a_528_n66# a_446_n108262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4975 a_2294_n80998# A1 a_2030_n80998# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4976 a_2030_n37688# A2 a_1634_n37688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4977 GND A5 word478 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4978 word880 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4979 GND A5 word67 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4980 word382 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4981 GND A8 word255 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4982 a_1370_n103008# a_1320_n66# a_1238_n103008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4983 a_2162_n122178# a_2112_n66# a_2030_n122178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4984 word733 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4985 GND A9 word471 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4986 GND A7 word108 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4987 a_446_n32860# A8 a_182_n32860# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4988 a_1766_n23346# A3 a_1502_n23346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4989 GND A1 word248 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4990 GND A9 word23 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4991 a_446_n79720# A8 a_50_n79720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4992 GND A7 word596 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4993 word885 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4994 GND A8 word252 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4995 a_1370_n102582# a_1320_n66# a_1238_n102582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X4996 a_2294_n126438# A1 a_2030_n126438# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4997 a_446_n18376# A8 a_182_n18376# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X4998 word874 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X4999 GND A7 word54 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5000 word815 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5001 GND A9 word190 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5002 GND A4 word803 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5003 GND A5 word706 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5004 GND A2 word313 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5005 a_2030_n75460# A2 a_1766_n75460# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5006 a_578_n137656# a_528_n66# a_314_n137656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5007 a_1502_n111244# A4 a_1238_n111244# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5008 GND A4 word744 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5009 word38 A0 a_2162_n5596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5010 word648 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5011 a_446_n87672# A8 a_50_n87672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5012 word589 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5013 word999 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5014 word855 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5015 a_1370_n13548# a_1320_n66# a_1238_n13548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5016 GND A7 word374 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5017 GND A5 word977 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5018 word940 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5019 GND A0 word784 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5020 word157 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5021 GND A7 word315 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5022 a_1238_n109256# A5 a_974_n109256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5023 a_1106_n8294# a_1056_n66# a_974_n8294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5024 word87 a_2376_n66# a_2162_n12554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5025 a_1766_n52740# A3 a_1370_n52740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5026 word871 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5027 GND A3 word947 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5028 a_1238_n131692# A5 a_974_n131692# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5029 word669 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5030 word947 a_2376_n66# a_2162_n134674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5031 word736 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5032 word753 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5033 GND A8 word577 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5034 word417 a_2376_n66# a_2294_n59414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5035 GND A8 word518 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5036 a_50_n108404# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5037 GND A0 word336 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5038 word719 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5039 a_1370_n140354# a_1320_n66# a_1238_n140354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5040 a_1766_n29878# A3 a_1370_n29878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5041 GND A7 word371 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5042 GND A9 word69 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5043 GND A2 word579 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5044 a_1238_n100168# A5 a_842_n100168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5045 GND A3 word725 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5046 a_578_n33712# a_528_n66# a_446_n33712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5047 GND A2 word88 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5048 GND A2 word147 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5049 a_1106_n41664# a_1056_n66# a_974_n41664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5050 word725 a_2376_n66# a_2294_n103150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5051 a_1370_n117492# a_1320_n66# a_1106_n117492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5052 word12 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5053 word979 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5054 a_1238_n138650# A5 a_842_n138650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5055 word353 a_2376_n66# a_2294_n50326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5056 word364 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5057 GND A2 word418 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5058 a_974_n72904# A6 a_710_n72904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5059 a_1106_n88524# a_1056_n66# a_842_n88524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5060 GND A4 word908 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5061 GND A7 word90 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5062 a_710_n114368# A7 a_314_n114368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5063 GND A1 word289 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5064 GND A2 word576 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5065 a_1766_n20790# A3 a_1370_n20790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5066 GND A8 word135 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5067 word985 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5068 a_1766_n76028# A3 a_1370_n76028# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5069 GND A1 word560 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5070 GND A7 word637 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5071 GND A1 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5072 word976 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5073 word783 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5074 a_446_n24198# A8 a_182_n24198# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5075 GND A1 word128 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5076 a_182_n23914# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5077 a_842_n89802# a_792_n66# a_710_n89802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5078 word1016 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5079 word915 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5080 GND A8 word682 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5081 GND A8 word623 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5082 GND A4 word844 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5083 GND A2 word354 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5084 word531 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5085 word822 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5086 a_578_n143478# a_528_n66# a_314_n143478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5087 a_710_n4318# A7 a_446_n4318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5088 GND A1 word616 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5089 a_2294_n109398# A1 a_2030_n109398# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5090 GND A3 word17 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5091 word54 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5092 a_446_n93494# A8 a_50_n93494# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5093 a_842_n11418# a_792_n66# a_710_n11418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5094 a_974_n18518# A6 a_578_n18518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5095 GND A2 word625 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5096 a_974_n40954# A6 a_710_n40954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5097 a_1370_n66230# a_1320_n66# a_1238_n66230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5098 word735 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5099 a_710_n3892# A7 a_446_n3892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5100 word399 a_2376_n66# a_2162_n56858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5101 a_50_n105848# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5102 a_50_n114226# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5103 GND A0 word436 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5104 word990 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5105 a_842_n10992# a_792_n66# a_710_n10992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5106 a_1766_n44078# A3 a_1370_n44078# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5107 a_1106_n25050# a_1056_n66# a_974_n25050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5108 word941 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5109 word888 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5110 a_182_n47202# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5111 a_1898_n21642# a_1848_n66# a_1766_n21642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5112 word306 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5113 a_182_n38824# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5114 word1020 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5115 GND A2 word459 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5116 GND A6 word641 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5117 GND A5 word852 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5118 a_182_n3608# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5119 GND A2 word400 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5120 a_1502_n123598# A4 a_1106_n123598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5121 a_710_n120190# A7 a_314_n120190# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5122 a_1370_n34280# a_1320_n66# a_1106_n34280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5123 GND A0 word930 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5124 a_842_n17950# a_792_n66# a_710_n17950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5125 word665 a_2376_n66# a_2294_n94630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5126 GND A7 word520 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5127 a_50_n143620# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5128 word233 a_2376_n66# a_2294_n33286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5129 word301 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5130 a_974_n55864# A6 a_578_n55864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5131 a_2030_n1620# A2 a_1634_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5132 word84 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5133 GND A6 word421 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5134 word882 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5135 a_314_n45214# a_264_n66# a_182_n45214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5136 a_1502_n20222# A4 a_1238_n20222# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5137 GND A0 word152 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5138 GND A1 word169 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5139 a_314_n36836# a_264_n66# a_182_n36836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5140 word631 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5141 GND A8 word664 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5142 a_50_n129136# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5143 word922 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5144 GND A0 word482 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5145 word572 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5146 word863 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5147 GND A1 word657 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5148 word716 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5149 word808 A0 a_2294_n114936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5150 a_1370_n89092# a_1320_n66# a_1106_n89092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5151 word348 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5152 a_182_n15252# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5153 word79 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5154 a_974_n24340# A6 a_578_n24340# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5155 a_1106_n62396# a_1056_n66# a_974_n62396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5156 word201 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5157 word795 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5158 word574 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5159 word793 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5160 GND A4 word355 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5161 a_50_n76738# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5162 a_50_n85116# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5163 word411 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5164 word567 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5165 a_974_n93636# A6 a_578_n93636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5166 GND A0 word260 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5167 word499 a_2376_n66# a_2162_n71058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5168 GND A7 word295 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5169 GND A6 word687 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5170 GND A2 word763 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5171 a_50_n111670# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5172 a_50_n120048# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5173 a_1898_n2330# a_1848_n66# a_1634_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5174 word76 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5175 word181 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5176 GND A2 word921 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5177 word56 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5178 GND A4 word194 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5179 a_1370_n49190# a_1320_n66# a_1238_n49190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5180 word284 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5181 a_842_n72052# a_792_n66# a_578_n72052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5182 a_974_n79152# A6 a_710_n79152# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5183 word765 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5184 word406 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5185 a_842_n103008# a_792_n66# a_578_n103008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5186 word189 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5187 GND A0 word316 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5188 a_182_n53024# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5189 a_1106_n118202# a_1056_n66# a_974_n118202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5190 a_182_n44646# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5191 word467 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5192 a_578_n92216# a_528_n66# a_446_n92216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5193 a_1898_n65946# a_1848_n66# a_1634_n65946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5194 word972 A0 a_2294_n138224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5195 GND A3 word581 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5196 word821 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5197 a_578_n22494# a_528_n66# a_446_n22494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5198 a_1238_n12412# A5 a_842_n12412# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5199 a_842_n102582# a_792_n66# a_578_n102582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5200 a_842_n32150# a_792_n66# a_578_n32150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5201 word125 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5202 a_974_n39250# A6 a_710_n39250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5203 word898 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5204 GND A2 word970 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5205 a_1766_n3040# A3 a_1370_n3040# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5206 a_1634_n51604# a_1584_n66# a_1502_n51604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5207 a_974_n61686# A6 a_578_n61686# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5208 GND A6 word521 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5209 word679 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5210 a_578_n69354# a_528_n66# a_314_n69354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5211 GND A4 word460 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5212 a_314_n51036# a_264_n66# a_182_n51036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5213 word864 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5214 a_314_n42658# a_264_n66# a_182_n42658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5215 a_1634_n101304# a_1584_n66# a_1502_n101304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5216 GND A4 word33 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5217 word545 a_2376_n66# a_2294_n77590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5218 a_50_n126580# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5219 a_1634_n28742# a_1584_n66# a_1502_n28742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5220 a_1502_n64526# A4 a_1238_n64526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5221 word51 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5222 a_314_n135810# a_264_n66# a_50_n135810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5223 GND A4 word516 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5224 word674 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5225 word389 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5226 a_182_n12696# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5227 a_182_n21074# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5228 a_1898_n118912# a_1848_n66# a_1766_n118912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5229 word242 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5230 word802 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5231 GND A3 word198 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5232 a_578_n60266# a_528_n66# a_314_n60266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5233 a_842_n140354# a_792_n66# a_578_n140354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5234 a_182_n59556# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5235 a_50_n82560# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5236 a_1898_n33996# a_1848_n66# a_1634_n33996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5237 GND A3 word356 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5238 a_314_n143762# a_264_n66# a_50_n143762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5239 GND A5 word136 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5240 word82 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5241 word281 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5242 a_578_n98748# a_528_n66# a_446_n98748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5243 GND A2 word745 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5244 word513 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5245 word732 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5246 a_1238_n18944# A5 a_974_n18944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5247 GND A4 word235 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5248 a_842_n47060# a_792_n66# a_710_n47060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5249 a_1238_n2330# A5 a_974_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5250 a_974_n76596# A6 a_710_n76596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5251 word447 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5252 a_182_n50468# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5253 a_314_n57568# a_264_n66# a_182_n57568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5254 a_1106_n124024# a_1056_n66# a_842_n124024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5255 GND A4 word133 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5256 a_1502_n32576# A4 a_1106_n32576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5257 a_314_n112238# a_264_n66# a_50_n112238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5258 word508 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5259 a_1106_n115646# a_1056_n66# a_974_n115646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5260 word287 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5261 word449 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5262 word122 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5263 GND A3 word405 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5264 GND A0 word628 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5265 GND A5 word72 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5266 a_1502_n79436# A4 a_1106_n79436# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5267 word659 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5268 word954 A0 a_2162_n135668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5269 GND A4 word621 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5270 a_2030_n104002# A2 a_1634_n104002# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5271 word939 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5272 GND A5 word343 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5273 a_578_n66798# a_528_n66# a_314_n66798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5274 a_1238_n56716# A5 a_974_n56716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5275 a_50_n97470# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5276 GND A9 word336 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5277 word246 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5278 a_974_n112664# A6 a_710_n112664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5279 word837 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5280 word327 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5281 GND A0 word564 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5282 a_1502_n70348# A4 a_1106_n70348# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5283 word559 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5284 word430 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5285 a_1898_n124734# a_1848_n66# a_1634_n124734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5286 GND A7 word862 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5287 a_182_n65378# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5288 GND A3 word180 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5289 a_1502_n47486# A4 a_1238_n47486# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5290 a_314_n127148# a_264_n66# a_50_n127148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5291 word788 A0 a_2294_n112096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5292 a_182_n57000# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5293 word456 A0 a_2294_n64952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5294 a_314_n118770# a_264_n66# a_50_n118770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5295 word269 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5296 word21 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5297 word105 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5298 word451 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5299 a_1898_n95056# a_1848_n66# a_1634_n95056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5300 a_710_n12838# A7 a_446_n12838# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5301 word714 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5302 word593 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5303 word453 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5304 GND A9 word111 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5305 a_1634_n72336# a_1584_n66# a_1370_n72336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5306 a_710_n90512# A7 a_446_n90512# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5307 a_182_n7300# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5308 word161 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5309 word234 A0 a_2162_n33428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5310 word762 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5311 a_314_n63390# a_264_n66# a_182_n63390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5312 a_1634_n122036# a_1584_n66# a_1370_n122036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5313 word170 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5314 a_1634_n113658# a_1584_n66# a_1370_n113658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5315 a_2162_n63532# a_2112_n66# a_1898_n63532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5316 a_1898_n101162# a_1848_n66# a_1766_n101162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5317 a_974_n127574# A6 a_578_n127574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5318 word163 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5319 a_1634_n49474# a_1584_n66# a_1370_n49474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5320 word104 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5321 GND A6 word784 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5322 word658 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5323 a_1898_n139644# a_1848_n66# a_1766_n139644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5324 a_710_n50610# A7 a_314_n50610# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5325 a_2030_n101446# A2 a_1634_n101446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5326 word226 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5327 GND A5 word384 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5328 word388 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5329 GND A9 word436 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5330 GND A9 word377 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5331 a_2030_n139928# A2 a_1634_n139928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5332 GND A3 word502 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5333 word228 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5334 a_2294_n61544# A1 a_2030_n61544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5335 a_1766_n130272# A3 a_1370_n130272# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5336 a_1634_n40386# a_1584_n66# a_1370_n40386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5337 word600 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5338 word819 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5339 word186 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5340 a_1238_n48054# A5 a_842_n48054# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5341 a_1238_n39676# A5 a_974_n39676# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5342 a_1898_n130556# a_1848_n66# a_1766_n130556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5343 a_446_n13406# A8 a_182_n13406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5344 word126 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5345 word370 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5346 word429 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5347 a_1634_n78868# a_1584_n66# a_1502_n78868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5348 a_182_n342# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5349 GND A9 word155 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5350 a_182_n71200# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5351 word207 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5352 word280 A0 a_2294_n39960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5353 a_1106_n136378# a_1056_n66# a_974_n136378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5354 a_1634_n128568# a_1584_n66# a_1502_n128568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5355 word275 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5356 a_2162_n78442# a_2112_n66# a_1898_n78442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5357 word654 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5358 a_2030_n130840# A2 a_1634_n130840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5359 a_446_n82702# A8 a_50_n82702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5360 a_1898_n107694# a_1848_n66# a_1766_n107694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5361 GND A5 word218 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5362 GND A5 word159 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5363 word426 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5364 a_1766_n137230# A3 a_1502_n137230# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5365 GND A3 word119 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5366 a_1238_n30588# A5 a_842_n30588# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5367 a_2030_n56006# A2 a_1634_n56006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5368 a_2030_n116356# A2 a_1766_n116356# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5369 word494 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5370 GND A9 word211 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5371 GND A9 word152 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5372 word575 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5373 a_2162_n123740# a_2112_n66# a_1898_n123740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5374 word744 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5375 GND A9 word482 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5376 a_2162_n38540# a_2112_n66# a_1898_n38540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5377 GND A8 word62 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5378 a_2294_n76454# A1 a_2030_n76454# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5379 word333 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5380 a_446_n100452# A8 a_50_n100452# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5381 a_974_n133396# A6 a_578_n133396# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5382 a_710_n73472# A7 a_446_n73472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5383 word473 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5384 word751 a_2376_n66# a_2162_n106842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5385 a_1502_n91080# A4 a_1238_n91080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5386 word1006 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5387 word955 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5388 word114 A0 a_2162_n16388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5389 a_1898_n145466# a_1848_n66# a_1634_n145466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5390 a_2162_n131692# a_2112_n66# a_1898_n131692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5391 word812 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5392 a_1370_n112522# a_1320_n66# a_1238_n112522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5393 a_446_n28316# A8 a_182_n28316# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5394 a_578_n100736# a_528_n66# a_446_n100736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5395 a_446_n19938# A8 a_182_n19938# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5396 a_2162_n46492# a_2112_n66# a_1898_n46492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5397 GND A9 word260 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5398 word602 A0 a_2162_n85684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5399 a_1766_n105280# A3 a_1502_n105280# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5400 word700 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5401 word1011 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5402 a_1106_n13832# a_1056_n66# a_842_n13832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5403 a_2030_n24056# A2 a_1634_n24056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5404 a_446_n97612# A8 a_50_n97612# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5405 word538 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5406 GND A5 word264 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5407 GND A5 word323 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5408 word1010 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5409 a_2294_n135952# A1 a_1898_n135952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5410 word725 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5411 a_446_n107410# A8 a_50_n107410# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5412 word599 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5413 word941 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5414 GND A9 word316 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5415 a_1634_n93068# a_1584_n66# a_1502_n93068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5416 GND A9 word257 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5417 word1017 a_2376_n66# a_2294_n144614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5418 a_446_n10850# A8 a_182_n10850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5419 GND A1 word93 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5420 GND A6 word29 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5421 a_2030_n93352# A2 a_1766_n93352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5422 a_2162_n138650# a_2112_n66# a_1898_n138650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5423 word380 A0 a_2294_n54160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5424 word908 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5425 GND A8 word717 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5426 a_1106_n142200# a_1056_n66# a_842_n142200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5427 word789 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5428 a_1766_n39818# A3 a_1370_n39818# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5429 GND A8 word97 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5430 GND A8 word156 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5431 a_1766_n70632# A3 a_1370_n70632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5432 a_446_n106984# A8 a_50_n106984# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5433 GND A1 word581 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5434 word309 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5435 a_710_n88382# A7 a_446_n88382# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5436 GND A6 word930 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5437 word250 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5438 a_1238_n110108# A5 a_974_n110108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5439 GND A6 word26 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5440 GND A2 word217 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5441 a_1106_n51604# a_1056_n66# a_842_n51604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5442 a_1238_n101730# A5 a_842_n101730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5443 GND A7 word783 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5444 a_2030_n122178# A2 a_1634_n122178# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5445 a_2030_n113800# A2 a_1766_n113800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5446 word493 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5447 GND A5 word530 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5448 a_1238_n83270# A5 a_842_n83270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5449 GND A6 word769 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5450 a_1502_n127716# A4 a_1238_n127716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5451 a_710_n124308# A7 a_314_n124308# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5452 a_710_n115930# A7 a_314_n115930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5453 GND A3 word851 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5454 a_1766_n30730# A3 a_1370_n30730# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5455 a_710_n48480# A7 a_314_n48480# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5456 GND A8 word44 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5457 word851 a_2376_n66# a_2162_n121042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5458 GND A8 word205 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5459 word1 a_2376_n66# a_2294_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5460 word332 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5461 a_2162_n106700# a_2112_n66# a_1898_n106700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5462 word988 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5463 a_446_n34138# A8 a_182_n34138# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5464 word794 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5465 a_974_n1052# A6 a_710_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5466 a_446_n25760# A8 a_182_n25760# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5467 a_1766_n16246# A3 a_1370_n16246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5468 a_1634_n99600# a_1584_n66# a_1370_n99600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5469 a_710_n123882# A7 a_314_n123882# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5470 GND A1 word25 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5471 GND A1 word356 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5472 GND A8 word693 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5473 GND A2 word424 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5474 GND A8 word763 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5475 GND A0 word956 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5476 word835 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5477 GND A8 word202 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5478 GND A7 word546 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5479 GND A7 word63 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5480 a_2294_n141774# A1 a_1898_n141774# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5481 GND A7 word888 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5482 word824 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5483 a_2030_n68360# A2 a_1766_n68360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5484 word539 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5485 GND A0 word734 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5486 word107 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5487 GND A7 word265 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5488 GND A7 word324 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5489 a_974_n8010# A6 a_710_n8010# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5490 a_1766_n45640# A3 a_1502_n45640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5491 GND A1 word405 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5492 GND A1 word952 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5493 GND A3 word897 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5494 word619 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5495 word821 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5496 word897 a_2376_n66# a_2294_n127574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5497 a_1370_n75744# a_1320_n66# a_1238_n75744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5498 GND A8 word527 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5499 word861 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5500 word958 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5501 GND A7 word321 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5502 GND A1 word461 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5503 a_974_n7584# A6 a_710_n7584# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5504 GND A2 word529 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5505 a_1106_n95908# a_1056_n66# a_974_n95908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5506 GND A5 word922 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5507 GND A5 word863 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5508 GND A4 word960 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5509 a_1502_n133538# A4 a_1106_n133538# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5510 a_1106_n34564# a_1056_n66# a_842_n34564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5511 a_578_n26612# a_528_n66# a_446_n26612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5512 a_1370_n44220# a_1320_n66# a_1106_n44220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5513 word314 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5514 GND A8 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5515 GND A7 word99 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5516 word303 a_2376_n66# a_2162_n43226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5517 a_1502_n119054# A4 a_1238_n119054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5518 GND A0 word222 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5519 GND A1 word180 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5520 GND A9 word14 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5521 a_1370_n43794# a_1320_n66# a_1106_n43794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5522 a_842_n35842# a_792_n66# a_578_n35842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5523 word733 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5524 GND A7 word587 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5525 GND A8 word745 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5526 a_2294_n125160# A1 a_2030_n125160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5527 a_1766_n91364# A3 a_1502_n91364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5528 a_1370_n99032# a_1320_n66# a_1106_n99032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5529 a_182_n16814# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5530 a_446_n17098# A8 a_182_n17098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5531 word151 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5532 a_1766_n82986# A3 a_1502_n82986# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5533 GND A7 word45 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5534 a_1106_n72336# a_1056_n66# a_842_n72336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5535 word865 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5536 GND A2 word304 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5537 GND A6 word427 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5538 a_1370_n139786# a_1320_n66# a_1238_n139786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5539 word831 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5540 a_578_n136378# a_528_n66# a_314_n136378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5541 word36 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5542 a_1502_n101588# A4 a_1238_n101588# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5543 a_578_n128000# a_528_n66# a_314_n128000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5544 a_446_n6874# A8 a_182_n6874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5545 word63 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5546 a_446_n86394# A8 a_50_n86394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5547 a_1370_n12270# a_1320_n66# a_1238_n12270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5548 GND A5 word968 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5549 a_974_n42232# A6 a_710_n42232# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5550 GND A7 word365 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5551 a_50_n121610# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5552 a_2162_n2898# a_2112_n66# a_2030_n2898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5553 GND A6 word266 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5554 a_1370_n59130# a_1320_n66# a_1238_n59130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5555 word478 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5556 a_1370_n81566# a_1320_n66# a_1106_n81566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5557 a_50_n107126# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5558 a_2294_n8862# A1 a_1898_n8862# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5559 word349 a_2376_n66# a_2294_n49758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5560 GND A0 word386 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5561 word940 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5562 GND A1 word344 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5563 word712 A0 a_2294_n101304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5564 a_1370_n130698# a_1320_n66# a_1238_n130698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5565 a_1370_n67082# a_1320_n66# a_1238_n67082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5566 GND A2 word570 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5567 a_578_n32434# a_528_n66# a_446_n32434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5568 a_1898_n14542# a_1848_n66# a_1766_n14542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5569 a_1766_n97896# A3 a_1370_n97896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5570 a_1766_n910# A3 a_1502_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5571 a_974_n80004# A6 a_710_n80004# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5572 a_1106_n87246# a_1056_n66# a_842_n87246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5573 GND A7 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5574 word285 a_2376_n66# a_2294_n40670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5575 GND A2 word409 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5576 a_1106_n78868# a_1056_n66# a_974_n78868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5577 GND A6 word532 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5578 GND A4 word840 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5579 a_710_n113090# A7 a_314_n113090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5580 word934 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5581 word993 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5582 GND A4 word98 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5583 word685 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5584 a_1370_n27180# a_1320_n66# a_1106_n27180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5585 word615 a_2376_n66# a_2162_n87530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5586 GND A0 word880 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5587 a_50_n136520# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5588 a_842_n50042# a_792_n66# a_710_n50042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5589 a_974_n57142# A6 a_578_n57142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5590 word183 a_2376_n66# a_2162_n26186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5591 GND A7 word569 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5592 GND A4 word586 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5593 a_182_n22636# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5594 a_182_n31014# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5595 a_314_n38114# a_264_n66# a_182_n38114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5596 GND A0 word102 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5597 GND A6 word310 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5598 a_842_n88524# a_792_n66# a_710_n88524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5599 GND A8 word614 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5600 a_578_n70206# a_528_n66# a_314_n70206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5601 a_1898_n52314# a_1848_n66# a_1634_n52314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5602 word671 a_2376_n66# a_2162_n95482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5603 a_578_n142200# a_528_n66# a_314_n142200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5604 a_710_n3040# A7 a_446_n3040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5605 a_50_n144472# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5606 a_578_n61828# a_528_n66# a_314_n61828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5607 a_1898_n43936# a_1848_n66# a_1766_n43936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5608 a_842_n141916# a_792_n66# a_578_n141916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5609 word758 A0 a_2162_n107836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5610 a_2030_n2472# A2 a_1766_n2472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5611 GND A2 word675 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5612 a_842_n10140# a_792_n66# a_710_n10140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5613 word743 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5614 word456 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5615 GND A2 word874 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5616 word524 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5617 a_50_n78016# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5618 a_1898_n29452# a_1848_n66# a_1634_n29452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5619 GND A6 word307 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5620 word517 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5621 GND A6 word696 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5622 a_314_n67508# a_264_n66# a_182_n67508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5623 a_50_n104570# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5624 a_974_n25192# A6 a_578_n25192# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5625 word131 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5626 GND A0 word368 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5627 a_182_n60408# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5628 GND A4 word203 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5629 a_1502_n42516# A4 a_1106_n42516# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5630 GND A4 word361 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5631 a_1898_n81708# a_1848_n66# a_1634_n81708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5632 GND A0 word698 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5633 a_2030_n9430# A2 a_1766_n9430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5634 word932 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5635 a_1898_n3182# a_1848_n66# a_1766_n3182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5636 a_1898_n20364# a_1848_n66# a_1634_n20364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5637 a_1502_n200# A4 a_1238_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5638 a_182_n37546# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5639 a_1502_n19654# A4 a_1238_n19654# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5640 a_1502_n28032# A4 a_1238_n28032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5641 GND A6 word415 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5642 word417 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5643 GND A2 word450 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5644 a_314_n121752# a_264_n66# a_50_n121752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5645 GND A6 word573 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5646 a_182_n2330# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5647 a_1898_n58846# a_1848_n66# a_1634_n58846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5648 word627 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5649 a_1502_n1762# A4 a_1238_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5650 GND A3 word531 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5651 GND A3 word54 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5652 word134 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5653 GND A2 word979 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5654 word351 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5655 GND A0 word634 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5656 word710 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5657 word292 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5658 a_1634_n44504# a_1584_n66# a_1370_n44504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5659 word629 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5660 word873 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5661 word814 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5662 GND A4 word42 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5663 a_1502_n10566# A4 a_1238_n10566# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5664 a_842_n85968# a_792_n66# a_710_n85968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5665 word622 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5666 word854 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5667 a_50_n119480# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5668 GND A0 word414 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5669 word563 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5670 GND A2 word976 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5671 word858 A0 a_2162_n122036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5672 a_182_n66940# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5673 a_314_n128710# a_264_n66# a_50_n128710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5674 word504 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5675 word339 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5676 word462 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5677 word280 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5678 GND A0 word22 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5679 word70 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5680 GND A6 word190 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5681 a_1898_n96618# a_1848_n66# a_1766_n96618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5682 word784 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5683 word497 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5684 GND A2 word915 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5685 word192 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5686 word565 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5687 a_1370_n2472# a_1320_n66# a_1238_n2472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5688 a_1898_n26896# a_1848_n66# a_1634_n26896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5689 a_1898_n35274# a_1848_n66# a_1766_n35274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5690 word402 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5691 a_842_n124876# a_792_n66# a_710_n124876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5692 a_50_n75460# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5693 GND A3 word306 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5694 GND A9 word181 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5695 a_314_n136662# a_264_n66# a_50_n136662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5696 a_974_n92358# A6 a_578_n92358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5697 a_1106_n99600# a_1056_n66# a_974_n99600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5698 word231 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5699 a_2294_n33712# A1 a_1898_n33712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5700 word91 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5701 GND A2 word754 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5702 GND A6 word678 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5703 a_1898_n111102# a_1848_n66# a_1634_n111102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5704 word397 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5705 GND A0 word680 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5706 word174 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5707 a_1502_n86820# A4 a_1106_n86820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5708 GND A3 word84 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5709 a_182_n43368# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5710 GND A4 word673 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5711 a_1106_n108546# a_1056_n66# a_842_n108546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5712 a_1634_n109114# a_1584_n66# a_1370_n109114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5713 a_182_n34990# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5714 word399 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5715 word458 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5716 word959 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5717 a_1238_n3182# A5 a_974_n3182# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5718 a_1898_n64668# a_1848_n66# a_1766_n64668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5719 word668 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5720 word904 A0 a_2294_n128568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5721 a_1238_n11134# A5 a_842_n11134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5722 word175 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5723 GND A0 word68 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5724 word889 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5725 a_578_n68076# a_528_n66# a_314_n68076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5726 word670 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5727 a_578_n59698# a_528_n66# a_314_n59698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5728 a_1238_n49616# A5 a_842_n49616# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5729 a_842_n139786# a_792_n66# a_578_n139786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5730 a_314_n41380# a_264_n66# a_182_n41380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5731 a_1634_n100026# a_1584_n66# a_1370_n100026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5732 a_2162_n41522# a_2112_n66# a_2030_n41522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5733 a_2294_n48622# A1 a_1898_n48622# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5734 word196 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5735 word604 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5736 a_974_n98890# A6 a_578_n98890# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5737 word663 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5738 GND A0 word514 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5739 word277 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5740 word42 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5741 a_1502_n54870# A4 a_1238_n54870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5742 a_1766_n100310# A3 a_1502_n100310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5743 word380 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5744 a_1634_n138508# a_1584_n66# a_1502_n138508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5745 word751 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5746 word503 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5747 word562 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5748 word665 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5749 a_1898_n126012# a_1848_n66# a_1766_n126012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5750 a_2030_n10708# A2 a_1634_n10708# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5751 word76 A0 a_2294_n10992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5752 word233 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5753 word71 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5754 a_1238_n40528# A5 a_974_n40528# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5755 word496 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5756 GND A7 word812 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5757 a_182_n49900# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5758 a_182_n58278# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5759 GND A3 word130 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5760 word406 A0 a_2162_n57852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5761 word505 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5762 GND A9 word281 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5763 GND A9 word222 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5764 a_314_n142484# a_264_n66# a_50_n142484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5765 a_710_n14116# A7 a_446_n14116# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5766 word73 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5767 word342 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5768 a_578_n97470# a_528_n66# a_446_n97470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5769 a_1898_n79578# a_1848_n66# a_1634_n79578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5770 GND A2 word795 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5771 word213 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5772 GND A3 word677 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5773 GND A6 word956 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5774 a_2162_n70916# a_2112_n66# a_2030_n70916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5775 word438 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5776 a_1634_n65236# a_1584_n66# a_1502_n65236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5777 a_710_n83412# A7 a_446_n83412# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5778 word543 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5779 a_974_n134958# A6 a_578_n134958# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5780 a_2294_n16672# A1 a_1898_n16672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5781 a_1634_n56858# a_1584_n66# a_1502_n56858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5782 word184 A0 a_2294_n26328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5783 word1017 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5784 a_314_n56290# a_264_n66# a_182_n56290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5785 a_1634_n106558# a_1584_n66# a_1502_n106558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5786 a_1106_n114368# a_1056_n66# a_974_n114368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5787 GND A2 word19 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5788 a_1106_n105990# a_1056_n66# a_842_n105990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5789 word440 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5790 word499 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5791 word113 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5792 a_1898_n70490# a_1848_n66# a_1634_n70490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5793 a_1502_n78158# A4 a_1106_n78158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5794 word672 A0 a_2294_n95624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5795 a_1502_n69780# A4 a_1106_n69780# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5796 word485 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5797 a_710_n43510# A7 a_314_n43510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5798 a_2030_n25618# A2 a_1766_n25618# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5799 GND A5 word393 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5800 word930 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5801 GND A5 word334 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5802 a_2162_n110108# a_2112_n66# a_1898_n110108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5803 a_1238_n55438# A5 a_974_n55438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5804 a_2162_n101730# a_2112_n66# a_2030_n101730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5805 GND A9 word386 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5806 GND A3 word452 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5807 word610 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5808 GND A9 word327 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5809 a_2162_n16530# a_2112_n66# a_2030_n16530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5810 word645 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5811 a_1634_n94630# a_1584_n66# a_1370_n94630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5812 a_2030_n94914# A2 a_1634_n94914# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5813 a_1766_n123172# A3 a_1502_n123172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5814 a_974_n111386# A6 a_710_n111386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5815 word769 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5816 a_1766_n114794# A3 a_1502_n114794# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5817 a_1634_n33286# a_1584_n66# a_1502_n33286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5818 a_710_n51462# A7 a_314_n51462# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5819 word259 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5820 word550 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5821 word136 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5822 a_2162_n94204# a_2112_n66# a_1898_n94204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5823 word851 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5824 GND A1 word981 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5825 GND A8 word167 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5826 a_2162_n85826# a_2112_n66# a_2030_n85826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5827 a_1898_n123456# a_1848_n66# a_1766_n123456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5828 GND A6 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5829 word379 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5830 a_2162_n24482# a_2112_n66# a_2030_n24482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5831 a_710_n89944# A7 a_446_n89944# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5832 word506 A0 a_2162_n72052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5833 GND A7 word794 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5834 GND A7 word853 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5835 GND A9 word105 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5836 a_182_n64100# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5837 a_2030_n132118# A2 a_1766_n132118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5838 a_446_n75602# A8 a_50_n75602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5839 word383 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5840 a_1238_n93210# A5 a_974_n93210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5841 a_710_n11560# A7 a_446_n11560# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5842 a_2294_n113942# A1 a_2030_n113942# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5843 word72 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5844 word376 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5845 a_2294_n92216# A1 a_2030_n92216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5846 GND A3 word659 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5847 GND A1 word917 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5848 a_2294_n83838# A1 a_1898_n83838# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5849 a_2030_n109256# A2 a_1766_n109256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5850 word786 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5851 GND A9 word161 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5852 GND A9 word102 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5853 a_2294_n22494# A1 a_1898_n22494# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5854 a_710_n80856# A7 a_446_n80856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5855 a_1634_n62680# a_1584_n66# a_1370_n62680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5856 a_2030_n62964# A2 a_1634_n62964# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5857 word525 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5858 GND A5 word656 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5859 a_2162_n125018# a_2112_n66# a_1898_n125018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5860 GND A5 word597 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5861 word753 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5862 a_1238_n92784# A5 a_974_n92784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5863 GND A7 word286 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5864 GND A1 word756 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5865 a_974_n2614# A6 a_710_n2614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5866 a_2162_n53876# a_2112_n66# a_2030_n53876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5867 GND A9 word43 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5868 a_1370_n47912# a_1320_n66# a_1238_n47912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5869 word905 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5870 GND A6 word775 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5871 a_578_n102014# a_528_n66# a_446_n102014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5872 a_2030_n100168# A2 a_1766_n100168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5873 a_1898_n138366# a_1848_n66# a_1634_n138366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5874 word762 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5875 word590 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5876 word552 A0 a_2294_n78584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5877 a_1502_n105706# A4 a_1106_n105706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5878 GND A9 word368 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5879 word58 A0 a_2162_n8436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5880 word961 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5881 a_2294_n51888# A1 a_1898_n51888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5882 word219 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5883 word359 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5884 word960 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5885 a_1238_n38398# A5 a_974_n38398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5886 GND A3 word967 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5887 word490 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5888 word891 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5889 GND A9 word207 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5890 a_446_n12128# A8 a_182_n12128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5891 word689 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5892 word967 a_2376_n66# a_2162_n137514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5893 a_2030_n77874# A2 a_1766_n77874# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5894 GND A8 a_264_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X5895 GND A7 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5896 word330 A0 a_2162_n47060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5897 GND A8 word106 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5898 word739 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5899 word1016 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5900 a_1370_n134816# a_1320_n66# a_1106_n134816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5901 a_1106_n135100# a_1056_n66# a_974_n135100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5902 a_1634_n127290# a_1584_n66# a_1370_n127290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5903 a_578_n131408# a_528_n66# a_314_n131408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5904 a_2162_n68786# a_2112_n66# a_2030_n68786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5905 a_446_n108262# A8 a_50_n108262# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5906 a_2162_n77164# a_2112_n66# a_1898_n77164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5907 a_446_n1904# A8 a_182_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5908 a_446_n81424# A8 a_50_n81424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5909 GND A5 word150 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5910 a_1106_n44504# a_1056_n66# a_974_n44504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5911 a_1238_n103008# A5 a_842_n103008# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5912 a_578_n108546# a_528_n66# a_446_n108546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5913 word695 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5914 a_2030_n115078# A2 a_1634_n115078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5915 word443 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5916 a_1238_n76170# A5 a_974_n76170# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5917 word688 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5918 a_578_n130982# a_528_n66# a_314_n130982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5919 word735 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5920 GND A5 word772 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5921 GND A7 word110 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5922 a_710_n117208# A7 a_314_n117208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5923 GND A9 word473 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5924 GND A9 word414 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5925 a_1766_n23630# A3 a_1502_n23630# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5926 a_1766_n32008# A3 a_1502_n32008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5927 a_2294_n66798# A1 a_1898_n66798# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5928 a_2294_n75176# A1 a_2030_n75176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5929 GND A3 word742 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5930 GND A1 word797 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5931 a_1238_n102582# A5 a_842_n102582# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5932 GND A9 word25 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5933 a_1370_n53734# a_1320_n66# a_1106_n53734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5934 a_1370_n62112# a_1320_n66# a_1106_n62112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5935 a_1898_n144188# a_1848_n66# a_1766_n144188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5936 word744 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5937 a_446_n27038# A8 a_182_n27038# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5938 a_1370_n102866# a_1320_n66# a_1238_n102866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5939 a_446_n18660# A8 a_182_n18660# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5940 a_710_n116782# A7 a_314_n116782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5941 word977 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5942 GND A5 word708 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5943 GND A2 word315 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5944 GND A0 word906 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5945 GND A4 word805 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5946 a_578_n137940# a_528_n66# a_314_n137940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5947 a_446_n96334# A8 a_50_n96334# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5948 a_1766_n78442# A3 a_1502_n78442# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5949 word40 A0 a_2294_n5880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5950 a_1370_n22210# a_1320_n66# a_1238_n22210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5951 a_446_n87956# A8 a_50_n87956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5952 word218 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5953 word159 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5954 a_1106_n59414# a_1056_n66# a_974_n59414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5955 a_1238_n109540# A5 a_974_n109540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5956 GND A7 word838 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5957 GND A3 word1008 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5958 a_1106_n8578# a_1056_n66# a_974_n8578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5959 word89 a_2376_n66# a_2294_n12838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5960 word932 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5961 GND A1 word1004 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5962 a_1238_n140354# A5 a_842_n140354# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5963 GND A3 word949 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5964 GND A1 word84 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5965 GND A2 word371 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5966 word949 a_2376_n66# a_2294_n134958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5967 a_710_n6732# A7 a_446_n6732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5968 GND A6 word20 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5969 word489 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5970 word755 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5971 a_1370_n30162# a_1320_n66# a_1238_n30162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5972 GND A7 word274 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5973 GND A8 word579 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5974 a_1370_n21784# a_1320_n66# a_1238_n21784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5975 GND A8 word147 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5976 a_1370_n140638# a_1320_n66# a_1238_n140638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5977 a_842_n13832# a_792_n66# a_710_n13832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5978 GND A8 word88 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5979 GND A1 word572 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5980 a_2294_n103150# A1 a_1898_n103150# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5981 word771 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5982 a_1370_n77022# a_1320_n66# a_1238_n77022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5983 a_1106_n50326# a_1056_n66# a_842_n50326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5984 word908 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5985 word752 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5986 a_1106_n41948# a_1056_n66# a_974_n41948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5987 GND A8 word576 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5988 a_1370_n126154# a_1320_n66# a_1106_n126154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5989 a_1370_n117776# a_1320_n66# a_1106_n117776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5990 GND A2 word90 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5991 GND A7 word271 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5992 a_578_n105990# a_528_n66# a_446_n105990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5993 a_1766_n46492# A3 a_1502_n46492# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5994 word425 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X5995 word355 a_2376_n66# a_2162_n50610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5996 a_1106_n88808# a_1056_n66# a_842_n88808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5997 GND A4 word910 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X5998 a_974_n20222# A6 a_578_n20222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X5999 a_710_n123030# A7 a_314_n123030# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6000 a_578_n19512# a_528_n66# a_446_n19512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6001 GND A8 word35 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6002 word783 a_2376_n66# a_2162_n111386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6003 word253 a_2376_n66# a_2294_n36126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6004 a_842_n51604# a_792_n66# a_710_n51604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6005 word264 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6006 a_974_n58704# A6 a_578_n58704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6007 GND A7 word639 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6008 word844 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6009 GND A0 word172 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6010 GND A1 word189 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6011 GND A4 word966 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6012 GND A4 word907 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6013 GND A8 word684 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6014 a_1370_n45072# a_1320_n66# a_1106_n45072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6015 word1018 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6016 GND A8 word625 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6017 GND A0 word1006 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6018 a_842_n28742# a_792_n66# a_578_n28742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6019 GND A7 word537 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6020 GND A8 word754 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6021 a_1766_n84264# A3 a_1370_n84264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6022 GND A1 word677 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6023 a_446_n93778# A8 a_50_n93778# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6024 a_1766_n75886# A3 a_1370_n75886# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6025 a_2294_n140496# A1 a_1898_n140496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6026 GND A6 word436 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6027 GND A2 word195 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6028 a_578_n129278# a_528_n66# a_314_n129278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6029 a_446_n8152# A8 a_182_n8152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6030 a_446_n79294# A8 a_50_n79294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6031 a_50_n114510# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6032 a_974_n26754# A6 a_578_n26754# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6033 GND A4 word431 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6034 GND A6 word155 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6035 a_842_n66514# a_792_n66# a_578_n66514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6036 word852 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6037 a_1898_n30304# a_1848_n66# a_1766_n30304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6038 word890 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6039 a_50_n122462# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6040 word308 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6041 GND A1 word452 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6042 GND A2 word520 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6043 GND A6 word643 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6044 GND A5 word854 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6045 word301 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6046 a_1502_n132260# A4 a_1106_n132260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6047 a_578_n25334# a_528_n66# a_446_n25334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6048 a_1106_n33286# a_1056_n66# a_842_n33286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6049 a_842_n105422# a_792_n66# a_578_n105422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6050 GND A6 word152 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6051 GND A6 word541 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6052 word235 a_2376_n66# a_2162_n33570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6053 a_1502_n109398# A4 a_1238_n109398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6054 word943 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6055 GND A4 word1007 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6056 word1019 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6057 word884 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6058 a_1502_n20506# A4 a_1238_n20506# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6059 GND A0 word830 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6060 a_50_n129420# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6061 a_842_n34564# a_792_n66# a_578_n34564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6062 GND A0 word484 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6063 GND A7 word578 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6064 GND A0 word988 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6065 a_1766_n5454# A3 a_1502_n5454# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6066 word47 a_2376_n66# a_2162_n6874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6067 word133 a_2376_n66# a_2294_n19086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6068 word574 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6069 GND A7 word519 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6070 a_182_n15536# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6071 word83 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6072 GND A6 word260 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6073 a_1370_n89376# a_1320_n66# a_1106_n89376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6074 word957 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6075 a_1106_n71058# a_1056_n66# a_842_n71058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6076 word3 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6077 a_578_n54728# a_528_n66# a_314_n54728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6078 a_578_n63106# a_528_n66# a_314_n63106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6079 a_1898_n45214# a_1848_n66# a_1634_n45214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6080 a_1106_n62680# a_1056_n66# a_974_n62680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6081 word621 a_2376_n66# a_2294_n88382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6082 a_578_n135100# a_528_n66# a_314_n135100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6083 word763 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6084 a_50_n137372# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6085 word413 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6086 word472 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6087 GND A1 word557 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6088 a_446_n5596# A8 a_182_n5596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6089 a_50_n128994# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6090 a_974_n93920# A6 a_578_n93920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6091 word406 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6092 GND A5 word900 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6093 GND A2 word824 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6094 GND A6 word257 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6095 GND A6 word316 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6096 word58 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6097 a_50_n93352# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6098 a_974_n79436# A6 a_710_n79436# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6099 a_1370_n80288# a_1320_n66# a_1106_n80288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6100 a_50_n84974# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6101 a_842_n63958# a_792_n66# a_578_n63958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6102 a_842_n72336# a_792_n66# a_578_n72336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6103 a_1634_n6164# a_1584_n66# a_1502_n6164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6104 a_2294_n7584# A1 a_1898_n7584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6105 GND A0 word318 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6106 a_182_n53308# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6107 a_182_n44930# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6108 a_842_n49474# a_792_n66# a_710_n49474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6109 a_1898_n74608# a_1848_n66# a_1634_n74608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6110 word974 A0 a_2162_n138508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6111 word970 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6112 a_578_n31156# a_528_n66# a_446_n31156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6113 a_578_n22778# a_528_n66# a_446_n22778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6114 a_1898_n13264# a_1848_n66# a_1634_n13264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6115 word247 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6116 a_842_n102866# a_792_n66# a_578_n102866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6117 GND A3 word151 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6118 word188 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6119 a_182_n52882# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6120 a_314_n59982# a_264_n66# a_182_n59982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6121 a_2294_n11702# A1 a_2030_n11702# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6122 a_974_n61970# A6 a_578_n61970# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6123 a_1106_n77590# a_1056_n66# a_974_n77590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6124 a_314_n114652# a_264_n66# a_50_n114652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6125 a_578_n69638# a_528_n66# a_314_n69638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6126 GND A6 word523 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6127 a_314_n51320# a_264_n66# a_182_n51320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6128 GND A3 word481 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6129 a_1766_n118912# A3 a_1502_n118912# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6130 a_974_n115504# A6 a_710_n115504# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6131 GND A0 word584 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6132 a_1502_n64810# A4 a_1238_n64810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6133 word956 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6134 word823 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6135 a_1766_n2898# A3 a_1370_n2898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6136 GND A4 word577 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6137 word764 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6138 a_182_n3182# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6139 a_182_n21358# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6140 word146 A0 a_2162_n20932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6141 a_842_n87246# a_792_n66# a_710_n87246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6142 GND A4 word518 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6143 a_1370_n95198# a_1320_n66# a_1238_n95198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6144 a_182_n12980# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6145 a_314_n50894# a_264_n66# a_182_n50894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6146 a_50_n99884# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6147 word244 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6148 word82 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6149 a_578_n60550# a_528_n66# a_314_n60550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6150 a_1898_n51036# a_1848_n66# a_1766_n51036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6151 a_842_n140638# a_792_n66# a_578_n140638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6152 a_182_n59840# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6153 a_182_n68218# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6154 a_50_n143194# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6155 GND A4 word416 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6156 a_1898_n89518# a_1848_n66# a_1766_n89518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6157 word506 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6158 word447 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6159 GND A2 word865 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6160 word734 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6161 a_1898_n28174# a_1848_n66# a_1766_n28174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6162 word515 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6163 a_842_n126154# a_792_n66# a_710_n126154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6164 a_1238_n27606# A5 a_842_n27606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6165 word40 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6166 GND A3 word256 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6167 word508 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6168 GND A9 word131 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6169 a_182_n67792# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6170 a_50_n90796# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6171 a_974_n76880# A6 a_710_n76880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6172 a_314_n129562# a_264_n66# a_50_n129562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6173 a_314_n66230# a_264_n66# a_182_n66230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6174 a_1502_n9572# A4 a_1238_n9572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6175 a_1502_n41238# A4 a_1106_n41238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6176 GND A0 word300 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6177 a_1106_n124308# a_1056_n66# a_842_n124308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6178 GND A4 word135 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6179 a_1502_n32860# A4 a_1106_n32860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6180 word571 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6181 a_1106_n115930# a_1056_n66# a_974_n115930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6182 GND A4 word352 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6183 word510 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6184 a_1898_n80430# a_1848_n66# a_1766_n80430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6185 GND A0 word630 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6186 GND A5 word74 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6187 word124 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6188 GND A4 word623 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6189 GND A4 word682 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6190 a_182_n27890# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6191 a_182_n36268# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6192 GND A3 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6193 a_1502_n18376# A4 a_1238_n18376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6194 word408 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6195 word246 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6196 a_314_n120474# a_264_n66# a_50_n120474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6197 a_1106_n123882# a_1056_n66# a_842_n123882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6198 word187 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6199 a_1898_n57568# a_1848_n66# a_1766_n57568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6200 GND A6 word564 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6201 a_1502_n87672# A4 a_1106_n87672# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6202 GND A6 word801 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6203 word248 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6204 word839 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6205 a_1634_n43226# a_1584_n66# a_1502_n43226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6206 word329 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6207 a_974_n112948# A6 a_710_n112948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6208 word620 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6209 word997 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6210 word862 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6211 a_1238_n64952# A5 a_842_n64952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6212 word613 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6213 a_842_n84690# a_792_n66# a_710_n84690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6214 GND A0 word464 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6215 a_1502_n56148# A4 a_1238_n56148# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6216 word676 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6217 word790 A0 a_2162_n112380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6218 a_1502_n47770# A4 a_1238_n47770# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6219 GND A4 word457 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6220 word330 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6221 word23 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6222 a_1898_n95340# a_1848_n66# a_1634_n95340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6223 word183 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6224 word775 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6225 word446 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6226 a_842_n123598# a_792_n66# a_710_n123598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6227 GND A9 word231 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6228 a_974_n91080# A6 a_578_n91080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6229 word455 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6230 GND A9 word172 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6231 a_1634_n72620# a_1584_n66# a_1370_n72620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6232 a_2030_n72904# A2 a_1766_n72904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6233 a_314_n135384# a_264_n66# a_50_n135384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6234 a_1766_n101162# A3 a_1502_n101162# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6235 GND A6 word669 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6236 word671 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6237 GND A5 word667 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6238 a_1634_n11276# a_1584_n66# a_1502_n11276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6239 word163 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6240 GND A3 word627 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6241 GND A6 word906 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6242 a_1634_n122320# a_1584_n66# a_1370_n122320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6243 a_1766_n139644# A3 a_1370_n139644# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6244 a_974_n136236# A6 a_578_n136236# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6245 a_974_n127858# A6 a_578_n127858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6246 word224 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6247 a_1634_n49758# a_1584_n66# a_1370_n49758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6248 a_710_n76312# A7 a_446_n76312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6249 word388 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6250 a_1634_n58136# a_1584_n66# a_1370_n58136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6251 word511 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6252 word165 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6253 word651 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6254 word967 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6255 a_314_n49190# a_264_n66# a_182_n49190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6256 word134 A0 a_2162_n19228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6257 a_2162_n134532# a_2112_n66# a_2030_n134532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6258 a_182_n42090# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6259 a_1502_n24198# A4 a_1106_n24198# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6260 word292 A0 a_2294_n41664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6261 a_1106_n107268# a_1056_n66# a_842_n107268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6262 a_2030_n101730# A2 a_1634_n101730# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6263 a_2162_n49332# a_2112_n66# a_2030_n49332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6264 word390 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6265 word950 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6266 a_1634_n121894# a_1584_n66# a_1370_n121894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6267 a_1898_n63390# a_1848_n66# a_1634_n63390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6268 GND A3 word563 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6269 word622 A0 a_2162_n88524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6270 word600 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6271 a_2294_n70206# A1 a_1898_n70206# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6272 word558 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6273 word69 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6274 word880 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6275 a_1766_n130556# A3 a_1370_n130556# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6276 a_2030_n18518# A2 a_1766_n18518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6277 word126 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6278 word230 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6279 word429 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6280 a_1634_n40670# a_1584_n66# a_1370_n40670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6281 a_1238_n48338# A5 a_842_n48338# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6282 word551 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6283 word70 A0 a_2162_n10140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6284 a_1238_n39960# A5 a_974_n39960# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6285 GND A3 word402 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6286 word654 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6287 GND A9 word277 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6288 a_2294_n38966# A1 a_2030_n38966# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6289 a_2162_n40244# a_2112_n66# a_2030_n40244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6290 a_2294_n47344# A1 a_1898_n47344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6291 a_2030_n87814# A2 a_1634_n87814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6292 a_710_n111812# A7 a_314_n111812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6293 a_1766_n107694# A3 a_1370_n107694# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6294 a_1766_n116072# A3 a_1370_n116072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6295 a_2162_n31866# a_2112_n66# a_1898_n31866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6296 a_182_n626# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6297 a_710_n44362# A7 a_314_n44362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6298 a_1370_n25902# a_1320_n66# a_1106_n25902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6299 word209 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6300 a_1106_n145040# a_1056_n66# a_842_n145040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6301 GND A8 word117 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6302 word742 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6303 word435 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6304 word494 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6305 a_1898_n107978# a_1848_n66# a_1766_n107978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6306 word616 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6307 a_446_n21642# A8 a_182_n21642# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6308 GND A5 word220 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6309 a_1634_n95482# a_1584_n66# a_1370_n95482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6310 GND A7 word803 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6311 GND A6 word46 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6312 word428 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6313 GND A9 word213 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6314 a_1634_n145182# a_1584_n66# a_1370_n145182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6315 a_578_n140922# a_528_n66# a_314_n140922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6316 a_1898_n78300# a_1848_n66# a_1766_n78300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6317 a_1238_n86110# A5 a_842_n86110# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6318 word145 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6319 GND A9 word484 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6320 GND A3 word609 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6321 GND A6 word947 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6322 word335 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6323 a_446_n100736# A8 a_50_n100736# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6324 a_974_n133680# A6 a_578_n133680# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6325 GND A1 word808 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6326 a_1238_n112522# A5 a_974_n112522# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6327 a_710_n73756# A7 a_446_n73756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6328 a_2030_n64242# A2 a_1766_n64242# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6329 word475 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6330 a_710_n82134# A7 a_446_n82134# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6331 a_2030_n55864# A2 a_1634_n55864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6332 GND A5 word606 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6333 word1008 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6334 a_2162_n109540# a_2112_n66# a_2030_n109540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6335 a_1238_n85684# A5 a_842_n85684# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6336 a_1238_n94062# A5 a_974_n94062# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6337 a_2162_n140354# a_2112_n66# a_2030_n140354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6338 word700 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6339 a_1370_n112806# a_1320_n66# a_1238_n112806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6340 a_2162_n55154# a_2112_n66# a_2030_n55154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6341 a_710_n126722# A7 a_314_n126722# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6342 a_1766_n41522# A3 a_1502_n41522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6343 GND A8 word61 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6344 word599 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6345 word604 A0 a_2294_n85968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6346 a_2162_n117492# a_2112_n66# a_2030_n117492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6347 a_2030_n24340# A2 a_1634_n24340# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6348 a_2294_n144614# A1 a_2030_n144614# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6349 GND A5 word325 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6350 GND A9 word318 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6351 GND A2 word441 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6352 GND A9 word259 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6353 GND A4 word931 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6354 word911 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6355 a_2294_n53166# A1 a_1898_n53166# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6356 a_2030_n93636# A2 a_1766_n93636# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6357 word309 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6358 word910 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6359 word127 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6360 a_1370_n31724# a_1320_n66# a_1238_n31724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6361 a_2030_n32292# A2 a_1766_n32292# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6362 a_1370_n40102# a_1320_n66# a_1238_n40102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6363 a_710_n50184# A7 a_314_n50184# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6364 GND A8 word158 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6365 GND A8 word217 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6366 a_2162_n84548# a_2112_n66# a_2030_n84548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6367 word841 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6368 GND A1 word972 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6369 GND A1 word913 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6370 a_1238_n127432# A5 a_974_n127432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6371 a_1766_n70916# A3 a_1370_n70916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6372 a_710_n88666# A7 a_446_n88666# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6373 GND A7 word844 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6374 word881 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6375 GND A7 word785 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6376 word966 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6377 word822 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6378 GND A2 word160 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6379 word438 A0 a_2162_n62396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6380 GND A7 word341 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6381 word907 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6382 GND A8 word646 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6383 a_446_n74324# A8 a_50_n74324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6384 GND A1 word481 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6385 GND A8 word716 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6386 word847 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6387 GND A6 word830 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6388 a_2294_n112664# A1 a_2030_n112664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6389 word47 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6390 GND A7 word16 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6391 GND A3 word853 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6392 GND A6 word181 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6393 a_2030_n39250# A2 a_1766_n39250# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6394 a_2294_n82560# A1 a_1898_n82560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6395 word777 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6396 word853 a_2376_n66# a_2294_n121326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6397 GND A1 word849 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6398 GND A2 word216 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6399 word393 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6400 GND A4 word706 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6401 word697 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6402 word3 a_2376_n66# a_2162_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6403 word334 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6404 a_2030_n61686# A2 a_1766_n61686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6405 GND A5 word588 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6406 GND A5 word647 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6407 word990 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6408 GND A2 word546 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6409 a_1766_n16530# A3 a_1370_n16530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6410 GND A9 word34 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6411 a_974_n1336# A6 a_710_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6412 a_2162_n99458# a_2112_n66# a_2030_n99458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6413 a_1370_n104144# a_1320_n66# a_1238_n104144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6414 GND A8 word765 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6415 word888 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6416 a_1898_n137088# a_1848_n66# a_1766_n137088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6417 a_1766_n94204# A3 a_1370_n94204# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6418 GND A7 word116 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6419 a_710_n109682# A7 a_314_n109682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6420 GND A7 word65 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6421 GND A1 word256 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6422 word633 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6423 GND A5 word717 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6424 a_446_n33996# A8 a_182_n33996# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6425 GND A2 word265 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6426 GND A7 word890 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6427 GND A9 word359 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6428 a_578_n139218# a_528_n66# a_314_n139218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6429 GND A9 word300 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6430 a_446_n9714# A8 a_182_n9714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6431 a_446_n89234# A8 a_50_n89234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6432 a_2294_n127574# A1 a_2030_n127574# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6433 word168 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6434 GND A5 word11 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6435 word109 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6436 a_2162_n90370# a_2112_n66# a_2030_n90370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6437 a_2294_n97470# A1 a_1898_n97470# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6438 word882 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6439 GND A1 word1013 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6440 a_2162_n5738# a_2112_n66# a_1898_n5738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6441 GND A3 word899 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6442 GND A4 word811 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6443 GND A2 word321 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6444 a_2030_n76596# A2 a_1634_n76596# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6445 a_1370_n84406# a_1320_n66# a_1238_n84406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6446 word899 a_2376_n66# a_2162_n127858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6447 a_578_n138792# a_528_n66# a_314_n138792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6448 GND A8 word529 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6449 word922 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6450 word1007 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6451 word863 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6452 a_578_n130130# a_528_n66# a_314_n130130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6453 a_50_n132402# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6454 GND A7 word382 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6455 GND A0 word792 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6456 a_446_n80146# A8 a_50_n80146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6457 a_1766_n62254# A3 a_1370_n62254# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6458 a_974_n7868# A6 a_710_n7868# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6459 GND A5 word924 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6460 word761 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6461 a_1106_n43226# a_1056_n66# a_974_n43226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6462 GND A6 word281 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6463 GND A2 word99 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6464 a_1106_n34848# a_1056_n66# a_842_n34848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6465 a_578_n107268# a_528_n66# a_446_n107268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6466 word1016 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6467 GND A8 word526 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6468 a_5404_164# A9 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X6469 a_1766_n39392# A3 a_1370_n39392# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6470 GND A8 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6471 a_2294_n2614# A1 a_2030_n2614# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6472 word16 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6473 word305 a_2376_n66# a_2294_n43510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6474 GND A9 word464 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6475 a_1502_n119338# A4 a_1238_n119338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6476 GND A2 word587 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6477 GND A5 word921 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6478 GND A1 word788 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6479 GND A2 word786 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6480 a_1502_n141774# A4 a_1106_n141774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6481 word733 a_2376_n66# a_2294_n104286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6482 a_1370_n52456# a_1320_n66# a_1106_n52456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6483 word203 a_2376_n66# a_2162_n29026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6484 GND A8 word245 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6485 GND A7 word589 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6486 GND A0 word122 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6487 word361 a_2376_n66# a_2294_n51462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6488 a_1766_n91648# A3 a_1502_n91648# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6489 word735 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6490 a_1238_n139786# A5 a_842_n139786# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6491 a_50_n100452# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6492 word153 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6493 word212 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6494 a_1370_n99316# a_1320_n66# a_1106_n99316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6495 GND A1 word297 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6496 a_1106_n72620# a_1056_n66# a_842_n72620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6497 word691 a_2376_n66# a_2162_n98322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6498 word702 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6499 a_578_n145040# a_528_n66# a_314_n145040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6500 a_1502_n110250# A4 a_1238_n110250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6501 word991 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6502 a_50_n138934# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6503 a_446_n86678# A8 a_50_n86678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6504 a_446_n95056# A8 a_50_n95056# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6505 a_1766_n68786# A3 a_1502_n68786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6506 GND A5 word970 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6507 a_974_n42516# A6 a_710_n42516# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6508 GND A6 word386 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6509 word923 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6510 GND A3 word999 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6511 a_1106_n7300# a_1056_n66# a_974_n7300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6512 a_1106_n80572# a_1056_n66# a_974_n80572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6513 word864 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6514 word999 a_2376_n66# a_2162_n142058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6515 a_1238_n130698# A5 a_974_n130698# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6516 a_1370_n90228# a_1320_n66# a_1106_n90228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6517 a_710_n5454# A7 a_446_n5454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6518 a_50_n94914# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6519 a_1370_n81850# a_1320_n66# a_1106_n81850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6520 GND A8 word570 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6521 word638 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6522 a_842_n12554# a_792_n66# a_710_n12554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6523 a_50_n107410# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6524 a_974_n19654# A6 a_578_n19654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6525 GND A2 word891 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6526 GND A3 word838 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6527 GND A7 word364 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6528 GND A4 word322 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6529 GND A1 word504 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6530 a_1370_n58988# a_1320_n66# a_1238_n58988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6531 a_1370_n67366# a_1320_n66# a_1238_n67366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6532 word840 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6533 a_578_n32718# a_528_n66# a_446_n32718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6534 a_1898_n14826# a_1848_n66# a_1766_n14826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6535 word317 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6536 word407 a_2376_n66# a_2162_n57994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6537 a_1370_n116498# a_1320_n66# a_1106_n116498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6538 a_50_n106984# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6539 a_50_n115362# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6540 a_182_n62822# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6541 a_314_n69922# a_264_n66# a_182_n69922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6542 a_1106_n87530# a_1056_n66# a_842_n87530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6543 a_1106_n26186# a_1056_n66# a_974_n26186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6544 GND A6 word161 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6545 GND A2 word569 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6546 a_974_n57426# A6 a_578_n57426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6547 word185 a_2376_n66# a_2294_n26470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6548 a_842_n50326# a_792_n66# a_710_n50326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6549 word969 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6550 word893 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6551 a_182_n4744# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6552 GND A0 word104 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6553 a_182_n22920# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6554 a_314_n60834# a_264_n66# a_182_n60834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6555 a_842_n88808# a_792_n66# a_710_n88808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6556 word1009 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6557 GND A8 word675 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6558 GND A4 word97 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6559 GND A0 word938 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6560 word874 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6561 word815 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6562 a_842_n27464# a_792_n66# a_578_n27464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6563 word673 a_2376_n66# a_2294_n95766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6564 word727 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6565 GND A7 word528 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6566 a_50_n144756# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6567 a_446_n92500# A8 a_50_n92500# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6568 GND A1 word609 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6569 GND A1 word668 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6570 a_2030_n2756# A2 a_1766_n2756# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6571 word92 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6572 GND A4 word486 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6573 a_1502_n82702# A4 a_1238_n82702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6574 a_182_n30872# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6575 a_314_n37972# a_264_n66# a_182_n37972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6576 a_578_n56006# a_528_n66# a_314_n56006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6577 word871 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6578 a_710_n2898# A7 a_446_n2898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6579 a_314_n139502# a_264_n66# a_50_n139502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6580 GND A5 word909 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6581 GND A6 word698 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6582 word87 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6583 a_974_n25476# A6 a_578_n25476# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6584 GND A0 word370 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6585 GND A4 word205 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6586 word801 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6587 word641 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6588 GND A4 word363 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6589 GND A4 word422 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6590 word582 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6591 a_50_n77874# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6592 a_50_n86252# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6593 a_842_n65236# a_792_n66# a_578_n65236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6594 word148 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6595 a_974_n94772# A6 a_578_n94772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6596 word934 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6597 GND A0 word268 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6598 word507 a_2376_n66# a_2162_n72194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6599 a_182_n37830# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6600 a_182_n46208# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6601 a_50_n121184# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6602 a_1898_n3466# a_1848_n66# a_1766_n3466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6603 a_1502_n28316# A4 a_1238_n28316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6604 GND A0 word426 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6605 GND A2 word771 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6606 a_1502_n19938# A4 a_1238_n19938# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6607 GND A4 word261 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6608 a_1502_n50752# A4 a_1106_n50752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6609 a_314_n130414# a_264_n66# a_50_n130414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6610 word979 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6611 a_1106_n133822# a_1056_n66# a_974_n133822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6612 GND A5 word845 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6613 GND A4 word202 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6614 GND A6 word575 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6615 word351 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6616 word292 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6617 word629 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6618 a_578_n24056# a_528_n66# a_446_n24056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6619 a_842_n104144# a_792_n66# a_578_n104144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6620 a_1502_n97612# A4 a_1106_n97612# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6621 word773 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6622 GND A3 word101 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6623 a_974_n63248# A6 a_578_n63248# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6624 a_182_n45782# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6625 word294 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6626 a_974_n54870# A6 a_578_n54870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6627 GND A6 word414 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6628 a_578_n93352# a_528_n66# a_446_n93352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6629 word875 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6630 a_314_n44220# a_264_n66# a_182_n44220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6631 GND A2 word707 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6632 GND A4 word44 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6633 a_1502_n10850# A4 a_1238_n10850# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6634 GND A0 word534 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6635 word915 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6636 a_1766_n484# A3 a_1502_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6637 a_842_n33286# a_792_n66# a_578_n33286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6638 word565 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6639 word860 A0 a_2294_n122320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6640 word62 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6641 GND A4 word527 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6642 word709 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6643 word906 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6644 word687 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6645 a_182_n14258# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6646 GND A7 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6647 a_314_n52172# a_264_n66# a_182_n52172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6648 GND A0 word24 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6649 word96 A0 a_2294_n13832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6650 word253 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6651 a_314_n43794# a_264_n66# a_182_n43794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6652 word91 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6653 word194 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6654 word754 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6655 a_1370_n2756# a_1320_n66# a_1238_n2756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6656 a_50_n136094# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6657 a_1898_n9998# a_1848_n66# a_1766_n9998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6658 word404 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6659 GND A3 word308 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6660 a_1502_n65662# A4 a_1238_n65662# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6661 a_314_n145324# a_264_n66# a_50_n145324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6662 word916 A0 a_2294_n130272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6663 word93 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6664 a_314_n136946# a_264_n66# a_50_n136946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6665 a_1766_n102724# A3 a_1370_n102724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6666 GND A6 word680 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6667 word397 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6668 VDD A8 a_264_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X6669 a_842_n119054# a_792_n66# a_710_n119054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6670 a_1634_n12838# a_1584_n66# a_1370_n12838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6671 a_50_n83696# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6672 a_50_n92074# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6673 a_842_n71058# a_792_n66# a_578_n71058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6674 a_974_n78158# A6 a_710_n78158# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6675 word581 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6676 a_2162_n12412# a_2112_n66# a_1898_n12412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6677 a_2294_n19512# A1 a_2030_n19512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6678 word399 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6679 a_1634_n90512# a_1584_n66# a_1370_n90512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6680 a_314_n59130# a_264_n66# a_182_n59130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6681 GND A0 word250 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6682 a_182_n52030# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6683 a_1502_n34138# A4 a_1106_n34138# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6684 word362 A0 a_2162_n51604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6685 a_578_n99884# a_528_n66# a_446_n99884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6686 a_1106_n108830# a_1056_n66# a_842_n108830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6687 word521 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6688 a_1106_n117208# a_1056_n66# a_974_n117208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6689 GND A4 word302 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6690 word460 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6691 a_1634_n140212# a_1584_n66# a_1370_n140212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6692 word298 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6693 a_1634_n131834# a_1584_n66# a_1370_n131834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6694 a_1238_n3466# A5 a_974_n3466# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6695 a_842_n48196# a_792_n66# a_710_n48196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6696 word670 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6697 word291 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6698 a_842_n101588# a_792_n66# a_578_n101588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6699 word814 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6700 a_182_n29168# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6701 a_578_n21500# a_528_n66# a_446_n21500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6702 a_1238_n11418# A5 a_842_n11418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6703 a_314_n67082# a_264_n66# a_182_n67082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6704 a_2294_n10424# A1 a_2030_n10424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6705 GND A3 word83 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6706 a_578_n68360# a_528_n66# a_314_n68360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6707 a_314_n113374# a_264_n66# a_50_n113374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6708 GND A6 word514 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6709 a_1634_n108972# a_1584_n66# a_1370_n108972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6710 a_1106_n116782# a_1056_n66# a_974_n116782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6711 GND A5 word512 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6712 a_1766_n126012# A3 a_1370_n126012# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6713 a_974_n114226# A6 a_710_n114226# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6714 a_1238_n10992# A5 a_842_n10992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6715 word198 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6716 a_1634_n36126# a_1584_n66# a_1370_n36126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6717 a_710_n45924# A7 a_314_n45924# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6718 a_710_n54302# A7 a_314_n54302# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6719 word279 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6720 word356 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6721 GND A2 word1019 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6722 word947 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6723 word1006 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6724 a_2162_n112522# a_2112_n66# a_1898_n112522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6725 a_182_n20080# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6726 a_1238_n57852# A5 a_974_n57852# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6727 a_1898_n117918# a_1848_n66# a_1634_n117918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6728 a_2162_n27322# a_2112_n66# a_1898_n27322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6729 word235 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6730 word795 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6731 word498 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6732 word445 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6733 word740 A0 a_2294_n105280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6734 word626 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6735 word403 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6736 word75 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6737 a_314_n142768# a_264_n66# a_50_n142768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6738 a_1898_n88240# a_1848_n66# a_1634_n88240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6739 word725 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6740 word438 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6741 GND A5 word129 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6742 word215 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6743 word133 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6744 a_1238_n9998# A5 a_842_n9998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6745 GND A3 word679 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6746 GND A5 word287 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6747 GND A9 word122 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6748 GND A3 word247 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6749 a_314_n128284# a_264_n66# a_50_n128284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6750 a_2030_n134532# A2 a_1766_n134532# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6751 a_2294_n25334# A1 a_2030_n25334# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6752 a_1634_n65520# a_1584_n66# a_1502_n65520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6753 word113 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6754 a_1898_n96192# a_1848_n66# a_1766_n96192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6755 a_2162_n141916# a_2112_n66# a_1898_n141916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6756 a_710_n13974# A7 a_446_n13974# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6757 word931 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6758 a_1106_n123030# a_1056_n66# a_842_n123030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6759 a_1634_n115220# a_1584_n66# a_1502_n115220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6760 a_2162_n56716# a_2112_n66# a_1898_n56716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6761 a_974_n129136# A6 a_578_n129136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6762 word115 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6763 word601 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6764 word461 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6765 word674 A0 a_2162_n95908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6766 word610 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6767 GND A4 word614 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6768 word242 A0 a_2162_n34564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6769 word178 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6770 word171 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6771 GND A3 word454 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6772 GND A3 word513 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6773 GND A9 word329 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6774 word981 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6775 a_2294_n54728# A1 a_2030_n54728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6776 GND A1 word712 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6777 GND A6 word792 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6778 a_1766_n123456# A3 a_1502_n123456# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6779 word379 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6780 word239 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6781 word666 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6782 a_974_n111670# A6 a_710_n111670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6783 word830 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6784 a_1634_n33570# a_1584_n66# a_1502_n33570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6785 a_710_n51746# A7 a_314_n51746# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6786 a_2030_n42232# A2 a_1634_n42232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6787 a_2030_n102582# A2 a_1766_n102582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6788 word988 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6789 GND A5 word392 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6790 GND A5 word451 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6791 word853 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6792 a_1898_n123740# a_1848_n66# a_1766_n123740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6793 GND A7 word81 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6794 word706 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6795 a_710_n37262# A7 a_314_n37262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6796 GND A7 word855 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6797 word508 A0 a_2294_n72336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6798 word977 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6799 word14 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6800 word917 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6801 a_1634_n88382# a_1584_n66# a_1502_n88382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6802 a_1898_n131692# a_1848_n66# a_1634_n131692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6803 a_446_n14542# A8 a_182_n14542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6804 word74 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6805 word378 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6806 word437 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6807 GND A3 word288 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6808 GND A9 word163 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6809 a_2030_n109540# A2 a_1766_n109540# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6810 a_2030_n80004# A2 a_1766_n80004# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6811 GND A9 word104 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6812 a_2030_n140354# A2 a_1634_n140354# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6813 a_1634_n138082# a_1584_n66# a_1502_n138082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6814 GND A5 word658 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6815 a_2030_n131976# A2 a_1766_n131976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6816 a_578_n133822# a_528_n66# a_314_n133822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6817 word755 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6818 word95 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6819 a_2294_n78016# A1 a_1898_n78016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6820 GND A6 word897 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6821 a_2162_n62538# a_2112_n66# a_1898_n62538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6822 a_2294_n69638# A1 a_2030_n69638# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6823 word344 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6824 a_446_n102014# A8 a_50_n102014# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6825 GND A1 word817 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6826 a_710_n75034# A7 a_446_n75034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6827 a_1766_n129988# A3 a_1370_n129988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6828 a_2030_n57142# A2 a_1766_n57142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6829 word502 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6830 a_2030_n117492# A2 a_1634_n117492# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6831 word583 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6832 a_1898_n138650# a_1848_n66# a_1634_n138650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6833 a_2162_n124876# a_2112_n66# a_1898_n124876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6834 word752 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6835 a_710_n119622# A7 a_314_n119622# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6836 word219 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6837 a_1766_n34422# A3 a_1370_n34422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6838 a_2162_n39676# a_2112_n66# a_1898_n39676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6839 word554 A0 a_2162_n78868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6840 GND A9 word429 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6841 GND A9 word370 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6842 word60 A0 a_2294_n8720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6843 a_2294_n60550# A1 a_2030_n60550# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6844 word963 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6845 GND A0 word50 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6846 a_2030_n17240# A2 a_1634_n17240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6847 word490 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6848 a_1766_n120900# A3 a_1370_n120900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6849 a_446_n29452# A8 a_182_n29452# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6850 GND A5 word275 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6851 a_578_n101872# a_528_n66# a_446_n101872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6852 a_1238_n47060# A5 a_842_n47060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6853 word483 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6854 GND A9 word268 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6855 a_2030_n86536# A2 a_1766_n86536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6856 GND A9 word426 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6857 GND A9 word209 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6858 a_2162_n30588# a_2112_n66# a_1898_n30588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6859 word119 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6860 a_2294_n37688# A1 a_2030_n37688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6861 a_710_n110534# A7 a_314_n110534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6862 a_1502_n113942# A4 a_1106_n113942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6863 a_710_n43084# A7 a_314_n43084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6864 a_2030_n25192# A2 a_1766_n25192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6865 GND A8 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6866 word667 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6867 word1018 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6868 word733 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6869 GND A0 word862 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6870 GND A8 word108 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6871 a_446_n81708# A8 a_50_n81708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6872 a_1766_n63816# A3 a_1502_n63816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6873 a_446_n108546# A8 a_50_n108546# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6874 a_1898_n106700# a_1848_n66# a_1634_n106700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6875 word607 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6876 a_446_n11986# A8 a_182_n11986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6877 a_446_n20364# A8 a_182_n20364# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6878 GND A1 word101 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6879 GND A6 word37 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6880 a_2162_n139786# a_2112_n66# a_1898_n139786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6881 word831 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6882 word388 A0 a_2294_n55296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6883 GND A8 word596 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6884 a_578_n108830# a_528_n66# a_446_n108830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6885 GND A9 word145 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6886 word797 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6887 GND A6 word938 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6888 GND A5 word991 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6889 GND A9 word475 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6890 GND A6 word131 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6891 GND A8 word55 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6892 a_1238_n111244# A5 a_974_n111244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6893 a_1766_n144188# A3 a_1370_n144188# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6894 GND A3 word803 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6895 a_1238_n102866# A5 a_842_n102866# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6896 word803 a_2376_n66# a_2162_n114226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6897 GND A5 word538 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6898 word999 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6899 word431 a_2376_n66# a_2162_n61402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6900 word442 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6901 a_2162_n130698# a_2112_n66# a_1898_n130698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6902 a_1370_n111528# a_1320_n66# a_1238_n111528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6903 a_1502_n128852# A4 a_1238_n128852# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6904 a_710_n125444# A7 a_314_n125444# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6905 GND A1 word308 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6906 a_2162_n45498# a_2112_n66# a_1898_n45498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6907 a_1370_n39534# a_1320_n66# a_1238_n39534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6908 GND A8 word52 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6909 word654 A0 a_2162_n93068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6910 word838 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6911 a_1766_n87104# A3 a_1502_n87104# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6912 a_446_n96618# A8 a_50_n96618# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6913 a_2294_n143336# A1 a_2030_n143336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6914 a_2294_n134958# A1 a_1898_n134958# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6915 word861 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6916 a_446_n35274# A8 a_182_n35274# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6917 a_446_n26896# A8 a_182_n26896# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6918 word220 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6919 GND A2 word274 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6920 GND A7 word840 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6921 GND A1 word33 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6922 a_1106_n90512# a_1056_n66# a_842_n90512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6923 GND A3 word1010 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6924 word934 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6925 word993 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6926 GND A8 word701 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6927 GND A9 word309 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6928 a_1238_n140638# A5 a_842_n140638# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6929 GND A2 word432 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6930 a_2030_n92358# A2 a_1634_n92358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6931 GND A9 word250 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6932 a_1370_n30446# a_1320_n66# a_1238_n30446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6933 GND A8 word710 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6934 GND A8 word90 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6935 GND A8 word149 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6936 word832 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6937 GND A1 word904 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6938 a_446_n105990# A8 a_50_n105990# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6939 word773 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6940 a_2030_n69496# A2 a_1634_n69496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6941 a_1370_n77306# a_1320_n66# a_1238_n77306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6942 a_710_n87388# A7 a_446_n87388# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6943 word606 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6944 GND A6 word19 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6945 GND A2 word210 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6946 a_1106_n50610# a_1056_n66# a_842_n50610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6947 GND A0 word742 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6948 word957 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6949 GND A8 word637 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6950 word910 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6951 a_1370_n126438# a_1320_n66# a_1106_n126438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6952 a_50_n125302# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6953 word477 a_2376_n66# a_2294_n67934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6954 GND A7 word273 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6955 GND A7 word332 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6956 a_974_n9146# A6 a_710_n9146# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6957 a_50_n116924# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6958 a_446_n73046# A8 a_50_n73046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6959 a_1766_n55154# A3 a_1502_n55154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6960 GND A1 word413 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6961 GND A1 word472 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6962 GND A8 word707 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6963 a_1106_n36126# a_1056_n66# a_842_n36126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6964 word700 A0 a_2294_n99600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6965 a_974_n20506# A6 a_578_n20506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6966 GND A7 word7 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6967 GND A6 word172 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6968 GND A3 word785 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6969 word907 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6970 word785 a_2376_n66# a_2294_n111670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6971 a_50_n72904# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6972 word255 a_2376_n66# a_2162_n36410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6973 GND A0 word174 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6974 GND A2 word537 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6975 GND A2 word736 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6976 a_1502_n143052# A4 a_1106_n143052# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6977 GND A4 word968 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6978 a_710_n122888# A7 a_314_n122888# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6979 GND A4 word167 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6980 a_1370_n45356# a_1320_n66# a_1106_n45356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6981 GND A0 word1008 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6982 GND A5 word66 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6983 GND A8 word254 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6984 GND A7 word598 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6985 word67 a_2376_n66# a_2162_n9714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6986 GND A8 word195 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6987 a_2162_n98180# a_2112_n66# a_2030_n98180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6988 GND A7 word539 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6989 GND A7 word107 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6990 word311 a_2376_n66# a_2162_n44362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6991 a_1766_n84548# A3 a_1370_n84548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6992 a_182_n40812# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X6993 a_314_n47912# a_264_n66# a_182_n47912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6994 GND A1 word188 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6995 a_446_n8436# A8 a_182_n8436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6996 a_446_n79578# A8 a_50_n79578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6997 GND A5 word979 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X6998 a_2294_n126296# A1 a_2030_n126296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X6999 GND A6 word277 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7000 word873 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7001 GND A1 word945 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7002 a_2162_n4460# a_2112_n66# a_1898_n4460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7003 word814 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7004 GND A4 word802 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7005 a_50_n87814# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7006 GND A8 word520 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7007 word854 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7008 a_1634_n9004# a_1584_n66# a_1370_n9004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7009 word577 a_2376_n66# a_2294_n82134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7010 word588 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7011 GND A5 word976 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7012 a_50_n131124# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7013 GND A7 word314 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7014 GND A7 word373 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7015 GND A1 word513 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7016 GND A2 word841 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7017 a_974_n6590# A6 a_710_n6590# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7018 a_50_n122746# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7019 GND A4 word331 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7020 a_1766_n52598# A3 a_1370_n52598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7021 GND A0 word496 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7022 word362 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7023 GND A5 word915 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7024 a_1106_n33570# a_1056_n66# a_842_n33570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7025 a_578_n25618# a_528_n66# a_446_n25618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7026 a_50_n108262# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7027 a_842_n105706# a_792_n66# a_578_n105706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7028 word1007 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7029 word208 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7030 a_182_n55722# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7031 GND A6 word543 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7032 a_2294_n1336# A1 a_2030_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7033 GND A2 word578 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7034 a_578_n94914# a_528_n66# a_446_n94914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7035 GND A2 word777 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7036 word11 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7037 word262 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7038 GND A0 word990 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7039 a_842_n34848# a_792_n66# a_578_n34848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7040 word135 a_2376_n66# a_2162_n19370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7041 a_1106_n88382# a_1056_n66# a_842_n88382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7042 GND A7 word580 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7043 word978 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7044 a_182_n6022# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7045 a_1766_n5738# A3 a_1502_n5738# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7046 a_1370_n98038# a_1320_n66# a_1106_n98038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7047 a_182_n15820# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7048 a_314_n62112# a_264_n66# a_182_n62112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7049 word144 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7050 GND A1 word288 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7051 a_1370_n89660# a_1320_n66# a_1106_n89660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7052 word942 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7053 word1001 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7054 a_314_n53734# a_264_n66# a_182_n53734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7055 GND A4 word106 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7056 word959 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7057 word623 a_2376_n66# a_2162_n88666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7058 GND A0 word888 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7059 a_50_n137656# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7060 word474 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7061 a_446_n5880# A8 a_182_n5880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7062 GND A1 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7063 a_2030_n4034# A2 a_1634_n4034# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7064 a_446_n85400# A8 a_50_n85400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7065 word986 A0 a_2162_n140212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7066 word467 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7067 a_974_n41238# A6 a_710_n41238# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7068 a_182_n23772# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7069 GND A6 word318 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7070 a_578_n71342# a_528_n66# a_314_n71342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7071 GND A6 word259 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7072 a_710_n4176# A7 a_446_n4176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7073 word60 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7074 a_578_n62964# a_528_n66# a_314_n62964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7075 a_50_n93636# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7076 GND A3 word16 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7077 a_842_n72620# a_792_n66# a_578_n72620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7078 a_974_n79720# A6 a_710_n79720# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7079 word766 A0 a_2162_n108972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7080 a_1634_n6448# a_1584_n66# a_1502_n6448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7081 GND A2 word683 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7082 a_842_n11276# a_792_n66# a_710_n11276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7083 a_974_n18376# A6 a_578_n18376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7084 GND A0 word320 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7085 word751 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7086 GND A2 word882 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7087 word532 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7088 word591 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7089 a_50_n79152# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7090 a_1370_n66088# a_1320_n66# a_1238_n66088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7091 a_842_n49758# a_792_n66# a_710_n49758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7092 word943 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7093 word457 a_2376_n66# a_2294_n65094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7094 word884 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7095 a_578_n31440# a_528_n66# a_446_n31440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7096 a_182_n39108# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7097 a_50_n114084# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7098 a_1898_n13548# a_1848_n66# a_1634_n13548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7099 GND A3 word212 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7100 word249 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7101 GND A0 word376 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7102 a_182_n61544# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7103 a_314_n68644# a_264_n66# a_182_n68644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7104 a_314_n123314# a_264_n66# a_50_n123314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7105 a_1106_n126722# a_1056_n66# a_842_n126722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7106 GND A5 word795 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7107 a_314_n114936# a_264_n66# a_50_n114936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7108 GND A6 word525 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7109 a_1898_n82844# a_1848_n66# a_1766_n82844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7110 GND A3 word65 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7111 a_182_n38682# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7112 a_1238_n20932# A5 a_974_n20932# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7113 word303 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7114 a_974_n56148# A6 a_578_n56148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7115 word244 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7116 word1017 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7117 a_314_n37120# a_264_n66# a_182_n37120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7118 GND A0 word154 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7119 GND A4 word579 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7120 word825 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7121 a_182_n3466# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7122 a_182_n30020# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7123 a_1898_n59982# a_1848_n66# a_1766_n59982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7124 a_842_n87530# a_792_n66# a_710_n87530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7125 word143 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7126 a_50_n143478# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7127 GND A0 word642 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7128 word718 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7129 word696 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7130 word810 A0 a_2162_n115220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7131 a_2030_n1478# A2 a_1634_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7132 GND A1 word600 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7133 GND A4 word418 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7134 word508 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7135 a_314_n36694# a_264_n66# a_182_n36694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7136 a_314_n45072# a_264_n66# a_182_n45072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7137 word203 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7138 GND A4 word576 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7139 word449 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7140 a_1370_n4034# a_1320_n66# a_1238_n4034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7141 a_842_n126438# a_792_n66# a_710_n126438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7142 a_1898_n28458# a_1848_n66# a_1766_n28458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7143 GND A6 word300 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7144 GND A3 word258 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7145 a_1898_n50894# a_1848_n66# a_1766_n50894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7146 word571 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7147 word866 A0 a_2162_n123172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7148 a_314_n129846# a_264_n66# a_50_n129846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7149 a_314_n138224# a_264_n66# a_50_n138224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7150 word510 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7151 word691 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7152 GND A6 word689 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7153 word347 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7154 word78 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7155 a_974_n24198# A6 a_578_n24198# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7156 a_1898_n97754# a_1848_n66# a_1634_n97754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7157 word851 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7158 word792 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7159 GND A2 word923 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7160 GND A2 word864 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7161 a_1502_n9856# A4 a_1238_n9856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7162 word573 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7163 GND A4 word354 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7164 a_50_n76596# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7165 word349 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7166 word566 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7167 a_1634_n83412# a_1584_n66# a_1502_n83412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7168 a_974_n93494# A6 a_578_n93494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7169 word925 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7170 a_1898_n2188# a_1848_n66# a_1634_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7171 GND A0 word200 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7172 GND A4 word684 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7173 a_182_n9998# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7174 GND A3 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7175 GND A2 word48 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7176 a_1502_n18660# A4 a_1238_n18660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7177 word312 A0 a_2294_n44504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7178 a_1634_n133112# a_1584_n66# a_1502_n133112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7179 word410 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7180 a_1106_n132544# a_1056_n66# a_974_n132544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7181 a_1634_n124734# a_1584_n66# a_1502_n124734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7182 a_314_n120758# a_264_n66# a_50_n120758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7183 word283 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7184 word823 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7185 GND A0 word688 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7186 word764 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7187 word241 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7188 a_1502_n87956# A4 a_1106_n87956# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7189 a_1502_n96334# A4 a_1106_n96334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7190 word285 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7191 GND A5 word462 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7192 word407 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7193 word466 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7194 a_578_n92074# a_528_n66# a_446_n92074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7195 a_1238_n73614# A5 a_974_n73614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7196 word615 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7197 GND A4 word35 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7198 a_2162_n34706# a_2112_n66# a_2030_n34706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7199 word183 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7200 a_1634_n29026# a_1584_n66# a_1502_n29026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7201 a_710_n47202# A7 a_314_n47202# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7202 a_710_n38824# A7 a_314_n38824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7203 word897 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7204 GND A2 word969 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7205 a_1634_n51462# a_1584_n66# a_1502_n51462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7206 word678 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7207 word762 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7208 word455 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7209 GND A4 word459 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7210 word185 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7211 a_1898_n141632# a_1848_n66# a_1766_n141632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7212 a_1634_n89944# a_1584_n66# a_1370_n89944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7213 word671 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7214 GND A3 word358 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7215 GND A9 word174 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7216 a_2294_n32718# A1 a_1898_n32718# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7217 word84 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7218 a_1502_n64384# A4 a_1238_n64384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7219 a_314_n135668# a_264_n66# a_50_n135668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7220 a_314_n144046# a_264_n66# a_50_n144046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7221 word388 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7222 word511 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7223 word673 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7224 a_2030_n11844# A2 a_1766_n11844# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7225 word165 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7226 GND A3 word629 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7227 a_1238_n19228# A5 a_974_n19228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7228 GND A3 word197 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7229 a_1238_n50042# A5 a_842_n50042# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7230 a_1898_n110108# a_1848_n66# a_1766_n110108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7231 word390 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7232 a_1634_n58420# a_1584_n66# a_1370_n58420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7233 a_2030_n127432# A2 a_1766_n127432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7234 word653 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7235 a_710_n15252# A7 a_446_n15252# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7236 a_1634_n80856# a_1584_n66# a_1370_n80856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7237 word221 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7238 word294 A0 a_2162_n41948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7239 a_1634_n108120# a_1584_n66# a_1370_n108120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7240 a_5404_164# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X7241 word230 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7242 a_1238_n2188# A5 a_974_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7243 word551 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7244 word624 A0 a_2294_n88808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7245 a_1238_n10140# A5 a_842_n10140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7246 GND A3 word565 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7247 word192 A0 a_2294_n27464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7248 a_314_n112096# a_264_n66# a_50_n112096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7249 word612 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7250 word553 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7251 word507 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7252 GND A5 word71 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7253 word121 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7254 a_2294_n56006# A1 a_2030_n56006# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7255 GND A3 word404 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7256 a_1502_n79294# A4 a_1106_n79294# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7257 GND A9 word279 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7258 GND A9 word496 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7259 a_1766_n116356# A3 a_1370_n116356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7260 a_710_n53024# A7 a_314_n53024# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7261 GND A8 word17 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7262 a_1766_n107978# A3 a_1370_n107978# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7263 a_182_n910# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7264 a_710_n44646# A7 a_314_n44646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7265 a_1634_n26470# a_1584_n66# a_1370_n26470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7266 a_2030_n26754# A2 a_1634_n26754# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7267 GND A5 word401 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7268 word938 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7269 word35 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7270 GND A5 word342 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7271 word744 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7272 a_1898_n125018# a_1848_n66# a_1634_n125018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7273 a_2162_n111244# a_2112_n66# a_1898_n111244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7274 a_1238_n56574# A5 a_974_n56574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7275 a_2162_n102866# a_2112_n66# a_2030_n102866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7276 a_1898_n116640# a_1848_n66# a_1766_n116640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7277 a_2162_n26044# a_2112_n66# a_1898_n26044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7278 word618 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7279 a_446_n30304# A8 a_182_n30304# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7280 a_1766_n12412# A3 a_1370_n12412# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7281 a_2162_n17666# a_2112_n66# a_2030_n17666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7282 a_446_n21926# A8 a_182_n21926# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7283 word458 A0 a_2162_n65236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7284 GND A7 word805 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7285 GND A9 word215 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7286 word867 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7287 word335 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7288 word394 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7289 a_314_n141490# a_264_n66# a_50_n141490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7290 GND A8 word736 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7291 a_1634_n145466# a_1584_n66# a_1370_n145466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7292 a_1106_n144898# a_1056_n66# a_842_n144898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7293 a_2162_n86962# a_2112_n66# a_2030_n86962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7294 a_1898_n124592# a_1848_n66# a_1634_n124592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7295 a_2294_n115504# A1 a_1898_n115504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7296 word67 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7297 GND A7 word36 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7298 GND A6 word949 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7299 GND A7 word861 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7300 GND A9 word113 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7301 a_1238_n112806# A5 a_974_n112806# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7302 a_2294_n24056# A1 a_2030_n24056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7303 a_710_n82418# A7 a_446_n82418# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7304 a_2030_n133254# A2 a_1634_n133254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7305 a_2294_n15678# A1 a_1898_n15678# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7306 word1010 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7307 a_1238_n94346# A5 a_974_n94346# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7308 word922 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7309 a_710_n12696# A7 a_446_n12696# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7310 a_1238_n85968# A5 a_842_n85968# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7311 a_2294_n93352# A1 a_2030_n93352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7312 a_1766_n41806# A3 a_1502_n41806# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7313 a_2294_n84974# A1 a_1898_n84974# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7314 word452 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7315 a_1634_n72194# a_1584_n66# a_1370_n72194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7316 a_710_n81992# A7 a_446_n81992# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7317 word533 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7318 a_2162_n126154# a_2112_n66# a_1898_n126154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7319 word761 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7320 a_1766_n18944# A3 a_1502_n18944# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7321 GND A9 word379 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7322 GND A9 word51 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7323 GND A9 word320 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7324 GND A6 word783 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7325 word913 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7326 a_1766_n113800# A3 a_1502_n113800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7327 a_710_n50468# A7 a_314_n50468# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7328 GND A5 word31 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7329 GND A8 word160 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7330 a_2162_n93210# a_2112_n66# a_1898_n93210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7331 word844 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7332 word287 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7333 word843 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7334 a_1238_n127716# A5 a_974_n127716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7335 GND A7 word72 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7336 a_710_n88950# A7 a_446_n88950# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7337 a_1502_n106842# A4 a_1106_n106842# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7338 GND A9 word376 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7339 GND A4 word772 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7340 word66 A0 a_2162_n9572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7341 GND A1 word153 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7342 GND A1 word212 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7343 a_1370_n17524# a_1320_n66# a_1106_n17524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7344 word617 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7345 GND A0 word812 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7346 word440 A0 a_2294_n62680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7347 GND A7 word343 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7348 word968 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7349 a_2162_n626# a_2112_n66# a_2030_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7350 a_446_n74608# A8 a_50_n74608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7351 word849 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7352 GND A8 word216 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7353 a_2294_n121326# A1 a_1898_n121326# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7354 a_446_n13264# A8 a_182_n13264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7355 word697 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7356 word369 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7357 GND A7 word18 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7358 word338 A0 a_2162_n48196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7359 word779 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7360 GND A8 word546 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7361 GND A9 word154 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7362 GND A9 word95 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7363 GND A3 word855 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7364 GND A4 word708 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7365 word747 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7366 a_1370_n135952# a_1320_n66# a_1106_n135952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7367 word855 a_2376_n66# a_2162_n121610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7368 a_578_n132544# a_528_n66# a_314_n132544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7369 a_2030_n61970# A2 a_1766_n61970# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7370 GND A5 word649 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7371 word699 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7372 word5 a_2376_n66# a_2294_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7373 GND A5 word590 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7374 GND A3 word550 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7375 a_1238_n91790# A5 a_974_n91790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7376 GND A3 word753 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7377 a_2162_n61260# a_2112_n66# a_1898_n61260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7378 a_2294_n68360# A1 a_2030_n68360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7379 a_1238_n104144# A5 a_842_n104144# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7380 GND A1 word749 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7381 a_1766_n137088# A3 a_1502_n137088# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7382 a_974_n1620# A6 a_710_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7383 word753 a_2376_n66# a_2294_n107126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7384 word633 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7385 word392 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7386 word890 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7387 word381 a_2376_n66# a_2294_n54302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7388 a_578_n101020# a_528_n66# a_446_n101020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7389 a_1370_n104428# a_1320_n66# a_1238_n104428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7390 GND A7 word118 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7391 GND A1 word317 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7392 a_710_n118344# A7 a_314_n118344# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7393 a_710_n109966# A7 a_314_n109966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7394 word635 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7395 GND A9 word33 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7396 a_1106_n14116# a_1056_n66# a_842_n14116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7397 word1013 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7398 a_446_n89518# A8 a_50_n89518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7399 word811 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7400 a_446_n28174# A8 a_182_n28174# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7401 word170 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7402 a_578_n100594# a_528_n66# a_446_n100594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7403 a_446_n19796# A8 a_182_n19796# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7404 word943 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7405 GND A3 word960 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7406 word884 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7407 GND A9 word200 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7408 GND A4 word872 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7409 GND A5 word716 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7410 GND A4 word813 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7411 word924 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7412 GND A8 word99 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7413 a_2162_n76170# a_2112_n66# a_1898_n76170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7414 word1009 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7415 a_1238_n119054# A5 a_842_n119054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7416 GND A0 word794 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7417 a_446_n80430# A8 a_50_n80430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7418 a_446_n107268# A8 a_50_n107268# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7419 GND A1 word524 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7420 word97 a_2376_n66# a_2294_n13974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7421 a_1766_n62538# A3 a_1370_n62538# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7422 GND A1 word92 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7423 GND A6 word28 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7424 a_1106_n43510# a_1056_n66# a_974_n43510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7425 word556 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7426 word763 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7427 GND A8 word587 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7428 word921 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7429 a_50_n109824# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7430 a_50_n118202# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7431 a_1766_n48054# A3 a_1370_n48054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7432 word1018 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7433 word786 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7434 a_1766_n39676# A3 a_1370_n39676# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7435 a_2294_n104286# A1 a_1898_n104286# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7436 word18 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7437 word69 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7438 GND A2 word648 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7439 a_1106_n51462# a_1056_n66# a_842_n51462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7440 a_1238_n101588# A5 a_842_n101588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7441 word735 a_2376_n66# a_2162_n104570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7442 a_1370_n52740# a_1320_n66# a_1106_n52740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7443 word205 a_2376_n66# a_2294_n29310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7444 word492 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7445 a_1106_n98322# a_1056_n66# a_974_n98322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7446 word363 a_2376_n66# a_2162_n51746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7447 a_1106_n89944# a_1056_n66# a_842_n89944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7448 GND A0 word124 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7449 a_710_n115788# A7 a_314_n115788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7450 word1012 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7451 a_1502_n127574# A4 a_1238_n127574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7452 a_710_n124166# A7 a_314_n124166# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7453 a_50_n100736# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7454 a_1766_n30588# A3 a_1370_n30588# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7455 word693 a_2376_n66# a_2294_n98606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7456 GND A7 word548 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7457 GND A0 word958 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7458 a_1370_n29878# a_1320_n66# a_1238_n29878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7459 GND A8 word204 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7460 word995 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7461 word261 a_2376_n66# a_2294_n37262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7462 a_446_n95340# A8 a_50_n95340# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7463 a_1766_n77448# A3 a_1502_n77448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7464 GND A1 word629 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7465 word112 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7466 a_2294_n133680# A1 a_1898_n133680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7467 GND A1 word197 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7468 a_182_n33712# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7469 GND A8 word692 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7470 a_1106_n80856# a_1056_n66# a_974_n80856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7471 word925 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7472 word891 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7473 a_2030_n91080# A2 a_1766_n91080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7474 a_578_n144898# a_528_n66# a_314_n144898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7475 a_710_n5738# A7 a_446_n5738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7476 word836 A0 a_2294_n118912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7477 a_974_n342# A6 a_710_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7478 a_974_n19938# A6 a_578_n19938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7479 a_1370_n20790# a_1320_n66# a_1238_n20790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7480 GND A8 word140 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7481 word823 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7482 a_842_n12838# a_792_n66# a_710_n12838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7483 GND A1 word565 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7484 a_1370_n76028# a_1320_n66# a_1238_n76028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7485 a_314_n40102# a_264_n66# a_182_n40102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7486 a_1370_n67650# a_1320_n66# a_1238_n67650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7487 a_842_n90512# a_792_n66# a_710_n90512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7488 word538 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7489 a_974_n97612# A6 a_578_n97612# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7490 a_1370_n125160# a_1320_n66# a_1106_n125160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7491 GND A7 word323 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7492 word527 a_2376_n66# a_2162_n75034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7493 GND A8 word569 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7494 a_50_n115646# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7495 a_50_n124024# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7496 GND A0 word446 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7497 GND A7 word264 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7498 GND A1 word404 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7499 word312 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7500 a_578_n18518# a_528_n66# a_446_n18518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7501 a_1106_n26470# a_1056_n66# a_974_n26470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7502 GND A6 word163 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7503 word957 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7504 a_182_n48622# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7505 a_50_n80004# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7506 a_842_n50610# a_792_n66# a_710_n50610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7507 a_974_n57710# A6 a_578_n57710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7508 GND A0 word224 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7509 GND A2 word528 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7510 a_1106_n95766# a_1056_n66# a_974_n95766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7511 GND A6 word651 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7512 a_1502_n133396# A4 a_1106_n133396# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7513 GND A4 word900 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7514 a_1370_n44078# a_1320_n66# a_1106_n44078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7515 a_1766_n7016# A3 a_1370_n7016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7516 a_842_n27748# a_792_n66# a_578_n27748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7517 a_842_n36126# a_792_n66# a_578_n36126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7518 a_1370_n35700# a_1320_n66# a_1106_n35700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7519 GND A8 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7520 GND A7 word530 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7521 GND A0 word940 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7522 word94 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7523 word951 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7524 a_314_n46634# a_264_n66# a_182_n46634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7525 a_314_n55012# a_264_n66# a_182_n55012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7526 GND A4 word646 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7527 word892 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7528 GND A6 word429 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7529 a_1106_n104712# a_1056_n66# a_842_n104712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7530 word431 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7531 GND A0 word838 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7532 a_446_n7158# A8 a_182_n7158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7533 a_446_n78300# A8 a_50_n78300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7534 word936 A0 a_2294_n133112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7535 a_1502_n68502# A4 a_1106_n68502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7536 word417 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7537 a_182_n16672# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7538 a_974_n25760# A6 a_578_n25760# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7539 word148 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7540 GND A2 word993 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7541 GND A6 word268 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7542 a_1106_n72194# a_1056_n66# a_842_n72194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7543 word862 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7544 word643 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7545 a_578_n55864# a_528_n66# a_314_n55864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7546 a_578_n64242# a_528_n66# a_314_n64242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7547 GND A4 word424 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7548 GND A6 word426 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7549 word771 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7550 a_50_n86536# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7551 a_842_n65520# a_792_n66# a_578_n65520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7552 word636 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7553 word710 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7554 GND A0 word270 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7555 word509 a_2376_n66# a_2294_n72478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7556 GND A2 word832 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7557 a_50_n121468# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7558 word541 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7559 GND A0 word428 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7560 GND A1 word445 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7561 GND A4 word263 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7562 word353 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7563 word294 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7564 word893 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7565 a_578_n24340# a_528_n66# a_446_n24340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7566 GND A6 word145 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7567 a_842_n104428# a_792_n66# a_578_n104428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7568 a_1766_n98180# A3 a_1370_n98180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7569 GND A0 word326 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7570 word707 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7571 a_182_n54444# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7572 GND A3 word103 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7573 GND A3 word162 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7574 a_1502_n36552# A4 a_1238_n36552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7575 a_314_n116214# a_264_n66# a_50_n116214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7576 GND A6 word534 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7577 a_1898_n84122# a_1848_n66# a_1634_n84122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7578 word477 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7579 GND A4 word1000 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7580 a_578_n93636# a_528_n66# a_446_n93636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7581 a_1898_n75744# a_1848_n66# a_1766_n75744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7582 a_578_n32292# a_528_n66# a_446_n32292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7583 word982 A0 a_2162_n139644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7584 word253 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7585 a_1766_n768# A3 a_1502_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7586 a_842_n33570# a_792_n66# a_578_n33570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7587 word967 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7588 a_1634_n61402# a_1584_n66# a_1502_n61402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7589 GND A7 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7590 word992 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7591 a_314_n52456# a_264_n66# a_182_n52456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7592 word933 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7593 word950 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7594 a_1634_n111102# a_1584_n66# a_1502_n111102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7595 word255 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7596 a_1898_n44220# a_1848_n66# a_1766_n44220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7597 word465 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7598 word760 A0 a_2294_n108120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7599 a_50_n128000# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7600 a_50_n136378# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7601 GND A0 word592 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7602 a_1502_n65946# A4 a_1238_n65946# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7603 a_1502_n74324# A4 a_1238_n74324# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7604 word918 A0 a_2162_n130556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7605 word458 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7606 word399 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7607 a_182_n22494# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7608 a_842_n88382# a_792_n66# a_710_n88382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7609 GND A4 word526 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7610 GND A6 word309 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7611 word252 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7612 a_842_n119338# a_792_n66# a_710_n119338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7613 a_578_n61686# a_528_n66# a_314_n61686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7614 a_578_n70064# a_528_n66# a_314_n70064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7615 a_1898_n52172# a_1848_n66# a_1634_n52172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7616 a_842_n141774# a_792_n66# a_578_n141774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7617 a_182_n69354# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7618 a_50_n92358# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7619 GND A3 word208 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7620 word460 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7621 word816 A0 a_2294_n116072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7622 a_50_n83980# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7623 GND A3 word7 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7624 a_2294_n6590# A1 a_1898_n6590# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7625 GND A2 word873 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7626 a_710_n16814# A7 a_446_n16814# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7627 word291 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7628 word742 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7629 word523 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7630 a_1238_n28742# A5 a_842_n28742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7631 word481 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7632 a_842_n48480# a_792_n66# a_710_n48480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7633 a_1238_n3750# A5 a_974_n3750# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7634 a_1898_n12270# a_1848_n66# a_1766_n12270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7635 word293 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7636 a_1634_n67934# a_1584_n66# a_1370_n67934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7637 word516 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7638 a_1634_n76312# a_1584_n66# a_1370_n76312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7639 word262 A0 a_2162_n37404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7640 word240 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7641 a_182_n60266# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7642 a_314_n67366# a_264_n66# a_182_n67366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7643 GND A3 word144 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7644 a_1502_n42374# A4 a_1106_n42374# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7645 a_314_n122036# a_264_n66# a_50_n122036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7646 a_1106_n125444# a_1056_n66# a_842_n125444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7647 a_182_n51888# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7648 a_314_n58988# a_264_n66# a_182_n58988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7649 word139 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7650 word198 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7651 a_1502_n33996# A4 a_1106_n33996# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7652 a_1898_n59130# a_1848_n66# a_1634_n59130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7653 a_314_n113658# a_264_n66# a_50_n113658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7654 a_1634_n117634# a_1584_n66# a_1370_n117634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7655 a_1502_n2046# A4 a_1238_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7656 GND A5 word141 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7657 word191 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7658 a_1898_n81566# a_1848_n66# a_1634_n81566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7659 word1019 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7660 GND A6 word812 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7661 a_2030_n9288# A2 a_1766_n9288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7662 GND A5 word82 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7663 word686 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7664 a_974_n114510# A6 a_710_n114510# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7665 a_1634_n36410# a_1584_n66# a_1370_n36410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7666 word416 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7667 word1008 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7668 GND A5 word412 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7669 word949 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7670 a_182_n2188# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7671 a_1238_n66514# A5 a_842_n66514# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7672 a_1898_n67082# a_1848_n66# a_1766_n67082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7673 word626 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7674 a_50_n98890# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7675 word75 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7676 word133 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7677 GND A2 word978 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7678 a_50_n142200# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7679 word628 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7680 a_1634_n35984# a_1584_n66# a_1370_n35984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7681 word499 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7682 word440 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7683 word135 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7684 word621 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7685 word980 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7686 a_1898_n27180# a_1848_n66# a_1634_n27180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7687 a_842_n125160# a_792_n66# a_710_n125160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7688 word345 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7689 GND A9 word124 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7690 a_182_n66798# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7691 a_314_n128568# a_264_n66# a_50_n128568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7692 word682 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7693 word338 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7694 a_2030_n13122# A2 a_1634_n13122# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7695 word115 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7696 a_1898_n96476# a_1848_n66# a_1766_n96476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7697 word783 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7698 a_1898_n103008# a_1848_n66# a_1766_n103008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7699 word564 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7700 a_974_n129420# A6 a_578_n129420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7701 word340 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7702 word463 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7703 word603 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7704 GND A4 word675 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7705 a_2162_n127716# a_2112_n66# a_2030_n127716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7706 word171 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7707 word244 A0 a_2294_n34848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7708 word239 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7709 a_1106_n122888# a_1056_n66# a_842_n122888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7710 a_974_n128994# A6 a_578_n128994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7711 word232 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7712 GND A3 word515 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7713 word173 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7714 a_1502_n86678# A4 a_1106_n86678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7715 a_1766_n132118# A3 a_1502_n132118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7716 GND A6 word794 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7717 a_1766_n123740# A3 a_1502_n123740# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7718 GND A2 word81 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7719 a_2030_n42516# A2 a_1634_n42516# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7720 a_578_n104712# a_528_n66# a_446_n104712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7721 a_2030_n102866# A2 a_1766_n102866# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7722 word457 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7723 GND A5 word453 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7724 word855 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7725 word990 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7726 a_1238_n63958# A5 a_842_n63958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7727 a_1766_n109256# A3 a_1502_n109256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7728 word708 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7729 GND A9 word446 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7730 a_2162_n33428# a_2112_n66# a_2030_n33428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7731 a_2294_n71342# A1 a_1898_n71342# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7732 a_710_n37546# A7 a_314_n37546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7733 a_2030_n19654# A2 a_1634_n19654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7734 word238 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7735 word437 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7736 word510 A0 a_2162_n72620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7737 word888 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7738 word669 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7739 word753 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7740 a_1238_n49474# A5 a_842_n49474# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7741 GND A4 word450 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7742 word78 A0 a_2162_n11276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7743 word627 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7744 a_446_n23204# A8 a_182_n23204# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7745 a_1634_n97044# a_1584_n66# a_1502_n97044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7746 a_446_n14826# A8 a_182_n14826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7747 word439 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7748 a_1634_n88666# a_1584_n66# a_1502_n88666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7749 word408 A0 a_2294_n58136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7750 GND A9 word224 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7751 GND A3 word290 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7752 word566 A0 a_2162_n80572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7753 GND A9 word165 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7754 a_1634_n138366# a_1584_n66# a_1502_n138366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7755 word817 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7756 a_2294_n31440# A1 a_1898_n31440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7757 a_2030_n71910# A2 a_1634_n71910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7758 a_314_n134390# a_264_n66# a_50_n134390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7759 a_1766_n100168# A3 a_1502_n100168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7760 word664 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7761 word502 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7762 GND A5 word660 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7763 a_2030_n10566# A2 a_1634_n10566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7764 GND A6 word958 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7765 GND A7 word811 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7766 GND A6 word899 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7767 GND A2 word186 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7768 a_1238_n40386# A5 a_974_n40386# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7769 a_1106_n4744# a_1056_n66# a_974_n4744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7770 a_710_n75318# A7 a_446_n75318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7771 a_2030_n57426# A2 a_1766_n57426# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7772 word504 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7773 GND A9 word221 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7774 word960 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7775 a_2162_n133538# a_2112_n66# a_2030_n133538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7776 word462 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7777 a_2162_n48338# a_2112_n66# a_2030_n48338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7778 GND A3 word676 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7779 a_710_n119906# A7 a_314_n119906# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7780 a_1766_n34706# A3 a_1370_n34706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7781 a_1634_n65094# a_1584_n66# a_1502_n65094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7782 word483 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7783 a_446_n101872# A8 a_50_n101872# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7784 a_710_n74892# A7 a_446_n74892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7785 a_1502_n92500# A4 a_1238_n92500# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7786 word1016 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7787 word119 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7788 a_446_n29736# A8 a_182_n29736# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7789 GND A1 word53 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7790 word544 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7791 GND A9 word270 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7792 a_2294_n46350# A1 a_1898_n46350# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7793 GND A5 word786 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7794 a_2030_n86820# A2 a_1766_n86820# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7795 a_710_n110818# A7 a_314_n110818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7796 GND A9 word428 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7797 a_710_n43368# A7 a_314_n43368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7798 GND A8 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7799 word607 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7800 a_2030_n25476# A2 a_1766_n25476# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7801 GND A5 word333 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7802 word237 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7803 word296 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7804 a_1238_n55296# A5 a_974_n55296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7805 GND A8 word110 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7806 a_2162_n101588# a_2112_n66# a_2030_n101588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7807 word735 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7808 word167 a_2376_n66# a_2162_n23914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7809 a_446_n108830# A8 a_50_n108830# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7810 a_2162_n16388# a_2112_n66# a_2030_n16388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7811 word609 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7812 GND A9 word326 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7813 a_446_n20648# A8 a_182_n20648# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7814 GND A6 word39 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7815 a_1634_n94488# a_1584_n66# a_1370_n94488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7816 a_2030_n94772# A2 a_1634_n94772# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7817 word390 A0 a_2162_n55580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7818 GND A0 word762 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7819 word991 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7820 word799 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7821 GND A8 word166 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7822 GND A8 word727 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7823 a_2162_n85684# a_2112_n66# a_2030_n85684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7824 a_2294_n105848# A1 a_2030_n105848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7825 word319 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7826 GND A7 word27 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7827 GND A7 word852 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7828 GND A6 word940 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7829 GND A1 word860 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7830 GND A3 word805 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7831 a_1238_n111528# A5 a_974_n111528# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7832 GND A2 word227 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7833 a_1106_n61402# a_1056_n66# a_974_n61402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7834 GND A4 word717 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7835 word805 a_2376_n66# a_2294_n114510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7836 a_2294_n14400# A1 a_1898_n14400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7837 a_2030_n54870# A2 a_1766_n54870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7838 a_710_n81140# A7 a_446_n81140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7839 GND A5 word599 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7840 GND A5 word540 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7841 a_1238_n84690# A5 a_842_n84690# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7842 a_1238_n93068# A5 a_974_n93068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7843 a_1502_n137514# A4 a_1238_n137514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7844 GND A1 word916 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7845 a_710_n125728# A7 a_314_n125728# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7846 GND A8 word54 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7847 a_2294_n83696# A1 a_1898_n83696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7848 GND A1 word857 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7849 a_1370_n39818# a_1320_n66# a_1238_n39818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7850 a_710_n49900# A7 a_314_n49900# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7851 word840 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7852 word861 a_2376_n66# a_2294_n122462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7853 word331 a_2376_n66# a_2162_n47202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7854 a_1370_n70632# a_1320_n66# a_1106_n70632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7855 a_2162_n116498# a_2112_n66# a_2030_n116498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7856 GND A7 word127 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7857 word922 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7858 word863 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7859 a_1766_n26044# A3 a_1370_n26044# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7860 a_446_n35558# A8 a_182_n35558# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7861 GND A1 word208 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7862 GND A9 word42 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7863 a_974_n2472# A6 a_710_n2472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7864 GND A2 word434 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7865 a_2294_n129136# A1 a_1898_n129136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7866 word761 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7867 a_1766_n86962# A3 a_1502_n86962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7868 GND A5 word22 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7869 word120 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7870 a_1370_n30730# a_1320_n66# a_1238_n30730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7871 a_2030_n31298# A2 a_1634_n31298# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7872 GND A8 word210 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7873 GND A1 word965 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7874 word834 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7875 word893 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7876 GND A2 word273 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7877 a_2030_n69780# A2 a_1634_n69780# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7878 a_1502_n105564# A4 a_1106_n105564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7879 GND A1 word144 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7880 a_1370_n16246# a_1320_n66# a_1106_n16246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7881 GND A0 word744 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7882 word959 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7883 GND A8 word639 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7884 GND A7 word334 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7885 word900 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7886 a_446_n73330# A8 a_50_n73330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7887 a_1766_n55438# A3 a_1502_n55438# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7888 GND A8 word709 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7889 GND A1 word1021 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7890 GND A3 word966 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7891 a_2294_n120048# A1 a_1898_n120048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7892 a_2162_n6874# a_2112_n66# a_1898_n6874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7893 a_2294_n111670# A1 a_2030_n111670# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7894 a_1370_n85542# a_1320_n66# a_1238_n85542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7895 word907 a_2376_n66# a_2162_n128994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7896 a_182_n11702# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7897 a_1106_n36410# a_1056_n66# a_842_n36410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7898 GND A7 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7899 GND A8 word537 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7900 GND A6 word174 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7901 word968 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7902 a_1370_n134674# a_1320_n66# a_1106_n134674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7903 GND A5 word640 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7904 a_578_n131266# a_528_n66# a_314_n131266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7905 word690 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7906 a_446_n1762# A8 a_182_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7907 word27 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7908 a_446_n81282# A8 a_50_n81282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7909 GND A2 word539 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7910 GND A1 word740 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7911 GND A4 word970 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7912 a_1106_n44362# a_1056_n66# a_974_n44362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7913 GND A2 word107 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7914 a_1106_n35984# a_1056_n66# a_842_n35984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7915 a_1370_n54018# a_1320_n66# a_1106_n54018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7916 word31 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7917 GND A5 word68 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7918 GND A0 word1010 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7919 word383 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7920 a_974_n75602# A6 a_710_n75602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7921 a_1370_n103150# a_1320_n66# a_1238_n103150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7922 a_50_n102014# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7923 word313 a_2376_n66# a_2294_n44646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7924 a_710_n117066# A7 a_314_n117066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7925 GND A5 word771 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7926 GND A7 word109 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7927 word979 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7928 a_1766_n23488# A3 a_1502_n23488# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7929 GND A1 word249 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7930 GND A0 word908 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7931 GND A5 word710 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7932 a_1370_n53592# a_1320_n66# a_1106_n53592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7933 word945 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7934 a_446_n8720# A8 a_182_n8720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7935 a_446_n88240# A8 a_50_n88240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7936 GND A7 word597 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7937 a_182_n26612# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7938 GND A6 word279 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7939 word976 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7940 word875 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7941 GND A4 word804 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7942 GND A5 word707 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7943 a_4612_164# A6 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X7944 a_710_n7016# A7 a_446_n7016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7945 a_578_n65804# a_528_n66# a_314_n65804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7946 GND A2 word314 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7947 a_578_n137798# a_528_n66# a_314_n137798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7948 a_1502_n111386# A4 a_1238_n111386# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7949 GND A4 word745 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7950 GND A3 word36 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7951 word46 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7952 a_446_n96192# A8 a_50_n96192# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7953 word649 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7954 word915 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7955 a_1370_n13690# a_1320_n66# a_1238_n13690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7956 a_1370_n22068# a_1320_n66# a_1238_n22068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7957 word579 a_2376_n66# a_2162_n82418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7958 word590 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7959 word1000 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7960 GND A0 word844 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7961 a_842_n14116# a_792_n66# a_710_n14116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7962 a_50_n131408# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7963 GND A7 word375 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7964 GND A2 word843 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7965 word147 a_2376_n66# a_2162_n21074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7966 a_974_n43652# A6 a_710_n43652# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7967 a_1106_n59272# a_1056_n66# a_974_n59272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7968 GND A0 word498 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7969 a_1238_n109398# A5 a_974_n109398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7970 word1007 a_2376_n66# a_2162_n143194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7971 word737 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7972 word754 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7973 word488 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7974 a_842_n83412# a_792_n66# a_710_n83412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7975 GND A8 word578 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7976 a_1370_n118060# a_1320_n66# a_1106_n118060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7977 GND A8 word519 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7978 a_1370_n140496# a_1320_n66# a_1238_n140496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7979 a_50_n108546# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7980 a_1634_n8862# a_1584_n66# a_1370_n8862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7981 GND A0 word396 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7982 a_50_n130982# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7983 word722 A0 a_2162_n102724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7984 word262 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7985 GND A2 word779 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7986 a_1106_n50184# a_1056_n66# a_842_n50184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7987 a_578_n33854# a_528_n66# a_446_n33854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7988 a_1898_n15962# a_1848_n66# a_1634_n15962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7989 a_974_n81424# A6 a_710_n81424# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X7990 a_1106_n88666# a_1056_n66# a_842_n88666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7991 a_1106_n97044# a_1056_n66# a_974_n97044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7992 word980 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7993 GND A2 word419 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7994 GND A4 word909 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7995 a_182_n6306# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7996 word1020 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7997 word1003 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X7998 GND A4 word108 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X7999 a_842_n29026# a_792_n66# a_578_n29026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8000 GND A0 word890 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8001 a_974_n58562# A6 a_578_n58562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8002 GND A1 word620 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8003 word625 a_2376_n66# a_2294_n88950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8004 GND A0 word662 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8005 a_50_n137940# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8006 a_842_n51462# a_792_n66# a_710_n51462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8007 a_1766_n76170# A3 a_1370_n76170# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8008 GND A7 word638 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8009 a_182_n32434# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8010 a_314_n39534# a_264_n66# a_182_n39534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8011 a_1502_n14542# A4 a_1106_n14542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8012 a_1370_n97896# a_1320_n66# a_1106_n97896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8013 a_842_n89944# a_792_n66# a_710_n89944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8014 GND A8 word683 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8015 a_1898_n62112# a_1848_n66# a_1766_n62112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8016 word882 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8017 GND A4 word845 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8018 a_578_n71626# a_528_n66# a_314_n71626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8019 word532 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8020 word886 A0 a_2162_n126012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8021 a_710_n4460# A7 a_446_n4460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8022 a_50_n93920# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8023 GND A1 word676 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8024 a_2030_n3892# A2 a_1634_n3892# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8025 GND A3 word18 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8026 a_974_n27038# A6 a_578_n27038# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8027 a_842_n11560# a_792_n66# a_710_n11560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8028 a_974_n18660# A6 a_578_n18660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8029 word812 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8030 a_578_n57142# a_528_n66# a_314_n57142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8031 word593 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8032 a_50_n79436# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8033 word795 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8034 GND A4 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8035 a_974_n96334# A6 a_578_n96334# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8036 word310 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8037 word459 a_2376_n66# a_2162_n65378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8038 a_182_n70206# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8039 a_50_n105990# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8040 a_50_n114368# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8041 GND A0 word378 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8042 a_182_n61828# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8043 a_314_n68928# a_264_n66# a_182_n68928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8044 a_1502_n52314# A4 a_1106_n52314# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8045 word303 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8046 GND A6 word154 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8047 a_842_n66372# a_792_n66# a_578_n66372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8048 word156 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8049 word942 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8050 GND A3 word112 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8051 GND A0 word276 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8052 a_182_n38966# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8053 a_182_n47344# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8054 a_1502_n29452# A4 a_1238_n29452# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8055 word307 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8056 word486 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8057 a_1898_n77022# a_1848_n66# a_1634_n77022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8058 word696 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8059 GND A6 word642 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8060 a_182_n3750# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8061 a_578_n25192# a_528_n66# a_446_n25192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8062 a_974_n132402# A6 a_578_n132402# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8063 word49 a_2376_n66# a_2294_n7158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8064 a_1634_n54302# a_1584_n66# a_1370_n54302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8065 GND A0 word644 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8066 word698 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8067 word85 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8068 GND A4 word420 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8069 word510 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8070 word883 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8071 a_314_n45356# a_264_n66# a_182_n45356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8072 a_1502_n20364# A4 a_1238_n20364# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8073 word205 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8074 a_1634_n104002# a_1584_n66# a_1370_n104002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8075 a_314_n36978# a_264_n66# a_182_n36978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8076 a_1898_n37120# a_1848_n66# a_1766_n37120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8077 word422 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8078 a_1370_n4318# a_1320_n66# a_1238_n4318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8079 a_50_n129278# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8080 word415 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8081 GND A0 word542 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8082 word923 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8083 word573 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8084 word868 A0 a_2294_n123456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8085 a_314_n138508# a_264_n66# a_50_n138508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8086 word693 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8087 word408 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8088 word531 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8089 word349 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8090 a_182_n15394# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8091 GND A0 word32 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8092 word853 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8093 word2 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8094 a_1898_n45072# a_1848_n66# a_1634_n45072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8095 word202 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8096 word575 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8097 word634 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8098 word794 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8099 a_842_n143052# a_792_n66# a_578_n143052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8100 a_1370_n3892# a_1320_n66# a_1238_n3892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8101 word471 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8102 a_50_n76880# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8103 a_50_n85258# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8104 a_974_n93778# A6 a_578_n93778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8105 word101 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8106 GND A6 word688 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8107 a_50_n120190# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8108 GND A3 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8109 a_1634_n22352# a_1584_n66# a_1370_n22352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8110 word241 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8111 a_1106_n141206# a_1056_n66# a_842_n141206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8112 word6 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8113 a_1106_n132828# a_1056_n66# a_974_n132828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8114 word57 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8115 GND A4 word195 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8116 word285 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8117 a_1898_n112522# a_1848_n66# a_1766_n112522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8118 a_842_n72194# a_792_n66# a_578_n72194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8119 a_974_n79294# A6 a_710_n79294# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8120 word243 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8121 word407 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8122 a_842_n103150# a_792_n66# a_578_n103150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8123 a_1502_n96618# A4 a_1106_n96618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8124 word190 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8125 a_182_n44788# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8126 a_182_n53166# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8127 a_2030_n112806# A2 a_1634_n112806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8128 word468 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8129 word306 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8130 a_578_n92358# a_528_n66# a_446_n92358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8131 GND A5 word91 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8132 GND A3 word641 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8133 GND A3 word582 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8134 word914 A0 a_2162_n129988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8135 a_1238_n12554# A5 a_842_n12554# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8136 word367 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8137 a_2294_n72904# A1 a_2030_n72904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8138 a_1766_n141632# A3 a_1502_n141632# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8139 a_1634_n29310# a_1584_n66# a_1502_n29310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8140 word958 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8141 word899 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8142 word55 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8143 a_1634_n51746# a_1584_n66# a_1502_n51746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8144 GND A4 word520 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8145 a_2162_n105706# a_2112_n66# a_1898_n105706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8146 word680 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8147 word148 A0 a_2294_n21216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8148 a_578_n69496# a_528_n66# a_314_n69496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8149 a_314_n42800# a_264_n66# a_182_n42800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8150 a_314_n51178# a_264_n66# a_182_n51178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8151 a_1634_n101446# a_1584_n66# a_1502_n101446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8152 a_1898_n141916# a_1848_n66# a_1766_n141916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8153 GND A3 word421 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8154 a_50_n135100# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8155 word206 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8156 a_974_n115362# A6 a_710_n115362# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8157 a_1634_n28884# a_1584_n66# a_1502_n28884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8158 a_1502_n73046# A4 a_1238_n73046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8159 a_1502_n64668# A4 a_1238_n64668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8160 a_314_n144330# a_264_n66# a_50_n144330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8161 word636 A0 a_2294_n90512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8162 a_1634_n139928# a_1584_n66# a_1370_n139928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8163 word850 A0 a_2162_n120900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8164 a_1766_n110108# A3 a_1502_n110108# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8165 a_2162_n89802# a_2112_n66# a_1898_n89802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8166 word390 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8167 a_842_n9714# a_792_n66# a_710_n9714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8168 a_182_n68076# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8169 GND A3 word199 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8170 GND A7 word822 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8171 GND A7 word881 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8172 a_842_n140496# a_792_n66# a_578_n140496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8173 a_182_n59698# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8174 a_50_n91080# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8175 a_2294_n18518# A1 a_2030_n18518# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8176 GND A9 word291 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8177 a_2030_n127716# A2 a_1766_n127716# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8178 a_2162_n11418# a_2112_n66# a_1898_n11418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8179 GND A3 word357 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8180 word411 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8181 a_710_n15536# A7 a_446_n15536# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8182 GND A2 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8183 a_578_n98890# a_528_n66# a_446_n98890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8184 a_1898_n89376# a_1848_n66# a_1766_n89376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8185 word733 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8186 GND A5 word137 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8187 word223 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8188 word83 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8189 GND A5 word196 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8190 word514 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8191 a_1238_n27464# A5 a_842_n27464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8192 GND A4 word295 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8193 a_1634_n130840# a_1584_n66# a_1370_n130840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8194 a_2162_n80714# a_2112_n66# a_1898_n80714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8195 a_2294_n87814# A1 a_2030_n87814# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8196 word472 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8197 a_1634_n75034# a_1584_n66# a_1502_n75034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8198 word553 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8199 a_710_n84832# A7 a_446_n84832# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8200 word121 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8201 word194 A0 a_2162_n27748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8202 a_314_n66088# a_264_n66# a_182_n66088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8203 a_1502_n41096# A4 a_1106_n41096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8204 a_1106_n124166# a_1056_n66# a_842_n124166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8205 a_1106_n115788# a_1056_n66# a_974_n115788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8206 word130 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8207 a_2162_n57852# a_2112_n66# a_1898_n57852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8208 a_314_n112380# a_264_n66# a_50_n112380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8209 word509 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8210 a_1898_n80288# a_1848_n66# a_1766_n80288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8211 GND A5 word73 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8212 word123 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8213 word182 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8214 GND A3 word465 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8215 word1014 A0 a_2162_n144188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8216 GND A6 word803 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8217 a_1502_n79578# A4 a_1106_n79578# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8218 GND A9 word498 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8219 a_1766_n116640# A3 a_1370_n116640# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8220 word618 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8221 a_710_n44930# A7 a_314_n44930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8222 a_2030_n35416# A2 a_1634_n35416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8223 a_710_n53308# A7 a_314_n53308# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8224 GND A5 word403 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8225 word940 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8226 word999 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8227 a_1238_n56858# A5 a_974_n56858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8228 a_1238_n65236# A5 a_842_n65236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8229 word611 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8230 word717 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8231 GND A9 word396 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8232 word247 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8233 word387 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8234 a_2294_n55864# A1 a_2030_n55864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8235 word838 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8236 a_710_n52882# A7 a_314_n52882# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8237 a_1634_n43084# a_1584_n66# a_1502_n43084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8238 word460 A0 a_2294_n65520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8239 word619 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8240 a_1502_n70490# A4 a_1106_n70490# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8241 GND A8 word236 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8242 word861 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8243 a_1898_n124876# a_1848_n66# a_1634_n124876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8244 a_446_n16104# A8 a_182_n16104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8245 GND A3 word240 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8246 GND A7 word863 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8247 GND A9 word115 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8248 word767 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8249 a_314_n127290# a_264_n66# a_50_n127290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8250 word516 A0 a_2294_n73472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8251 a_2030_n133538# A2 a_1634_n133538# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8252 word22 A0 a_2162_n3324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8253 a_1238_n94630# A5 a_974_n94630# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8254 a_1898_n95198# a_1848_n66# a_1634_n95198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8255 GND A6 word908 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8256 a_710_n12980# A7 a_446_n12980# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8257 word924 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8258 word141 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8259 a_1106_n6022# a_1056_n66# a_974_n6022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8260 GND A2 word136 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8261 word454 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8262 GND A9 word171 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8263 GND A3 word931 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8264 word931 a_2376_n66# a_2162_n132402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8265 word412 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8266 a_1634_n72478# a_1584_n66# a_1370_n72478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8267 a_710_n90654# A7 a_446_n90654# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8268 GND A5 word666 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8269 word763 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8270 GND A3 word626 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8271 word703 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8272 word921 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8273 a_1634_n122178# a_1584_n66# a_1370_n122178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8274 a_1766_n27606# A3 a_1502_n27606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8275 a_2162_n63674# a_2112_n66# a_1898_n63674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8276 a_2162_n72052# a_2112_n66# a_2030_n72052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8277 a_2294_n79152# A1 a_1898_n79152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8278 a_974_n136094# A6 a_578_n136094# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8279 GND A9 word53 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8280 word164 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8281 GND A6 word785 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8282 GND A1 word705 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8283 word966 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8284 word831 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8285 GND A2 word72 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8286 a_578_n103434# a_528_n66# a_446_n103434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8287 word659 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8288 a_1898_n139786# a_1848_n66# a_1766_n139786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8289 a_2030_n41238# A2 a_1766_n41238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8290 a_2030_n101588# A2 a_1634_n101588# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8291 GND A5 word385 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8292 GND A7 word74 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8293 a_2030_n79720# A2 a_1766_n79720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8294 GND A9 word437 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8295 GND A9 word378 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8296 a_1502_n115504# A4 a_1106_n115504# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8297 word68 A0 a_2294_n9856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8298 a_2294_n61686# A1 a_2030_n61686# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8299 a_2294_n70064# A1 a_1898_n70064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8300 GND A3 word706 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8301 a_2030_n18376# A2 a_1766_n18376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8302 a_1370_n17808# a_1320_n66# a_1106_n17808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8303 word369 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8304 a_2162_n79010# a_2112_n66# a_2030_n79010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8305 word970 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8306 word187 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8307 a_1238_n48196# A5 a_842_n48196# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8308 word117 a_2376_n66# a_2294_n16814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8309 GND A9 word276 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8310 GND A3 word977 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8311 a_1898_n130698# a_1848_n66# a_1766_n130698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8312 GND A1 word112 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8313 GND A6 word48 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8314 word430 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8315 word699 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8316 word977 a_2376_n66# a_2294_n138934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8317 a_446_n13548# A8 a_182_n13548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8318 a_2030_n87672# A2 a_1634_n87672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8319 a_182_n484# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8320 word340 A0 a_2294_n48480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8321 word749 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8322 a_1370_n144614# a_1320_n66# a_1106_n144614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8323 a_578_n141206# a_528_n66# a_314_n141206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8324 a_578_n132828# a_528_n66# a_314_n132828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8325 GND A8 word116 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8326 a_446_n91222# A8 a_50_n91222# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8327 a_2294_n107126# A1 a_2030_n107126# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8328 a_446_n82844# A8 a_50_n82844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8329 GND A5 word219 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8330 a_1106_n54302# a_1056_n66# a_842_n54302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8331 a_446_n101020# A8 a_50_n101020# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8332 a_1238_n104428# A5 a_842_n104428# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8333 GND A7 word802 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8334 GND A3 word755 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8335 GND A2 word177 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8336 a_710_n74040# A7 a_446_n74040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8337 a_2030_n56148# A2 a_1634_n56148# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8338 word495 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8339 word755 a_2376_n66# a_2162_n107410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8340 a_2030_n116498# A2 a_1766_n116498# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8341 word635 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8342 a_2162_n132260# a_2112_n66# a_2030_n132260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8343 GND A5 word841 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8344 a_2162_n47060# a_2112_n66# a_2030_n47060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8345 word745 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8346 GND A9 word483 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8347 a_710_n127006# A7 a_314_n127006# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8348 a_710_n118628# A7 a_314_n118628# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8349 GND A8 word63 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8350 a_446_n100594# A8 a_50_n100594# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8351 word811 a_2376_n66# a_2162_n115362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8352 GND A3 word752 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8353 a_1370_n63532# a_1320_n66# a_1106_n63532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8354 word1015 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8355 word1007 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8356 word872 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8357 a_2294_n136520# A1 a_2030_n136520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8358 a_1370_n121042# a_1320_n66# a_1238_n121042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8359 word813 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8360 a_1370_n112664# a_1320_n66# a_1238_n112664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8361 a_446_n28458# A8 a_182_n28458# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8362 a_578_n100878# a_528_n66# a_446_n100878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8363 GND A1 word44 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8364 GND A2 word443 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8365 GND A4 word874 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8366 GND A5 word777 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8367 GND A2 word384 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8368 GND A4 word815 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8369 a_1106_n13974# a_1056_n66# a_842_n13974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8370 a_710_n42090# A7 a_314_n42090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8371 a_2030_n24198# A2 a_1634_n24198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8372 a_446_n97754# A8 a_50_n97754# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8373 a_1766_n79862# A3 a_1370_n79862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8374 a_2294_n144472# A1 a_2030_n144472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8375 word217 a_2376_n66# a_2294_n31014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8376 a_1106_n69212# a_1056_n66# a_842_n69212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8377 a_1238_n119338# A5 a_842_n119338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8378 word600 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8379 word942 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8380 word1001 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8381 a_2030_n93494# A2 a_1766_n93494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8382 GND A4 word871 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8383 word824 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8384 GND A6 word30 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8385 word558 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8386 GND A8 word648 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8387 word765 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8388 word909 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8389 GND A8 word589 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8390 word126 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8391 a_1370_n31582# a_1320_n66# a_1238_n31582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8392 GND A8 word718 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8393 a_50_n140922# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8394 a_1766_n48338# A3 a_1370_n48338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8395 GND A8 word157 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8396 GND A1 word641 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8397 word49 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8398 a_1766_n70774# A3 a_1370_n70774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8399 a_1106_n60124# a_1056_n66# a_974_n60124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8400 a_1238_n110250# A5 a_974_n110250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8401 word821 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8402 GND A2 word218 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8403 a_1106_n51746# a_1056_n66# a_842_n51746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8404 a_1898_n25902# a_1848_n66# a_1766_n25902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8405 word336 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8406 a_446_n74182# A8 a_50_n74182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8407 GND A1 word421 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8408 word494 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8409 GND A2 word489 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8410 a_1106_n98606# a_1056_n66# a_974_n98606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8411 a_1502_n127858# A4 a_1238_n127858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8412 a_710_n124450# A7 a_314_n124450# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8413 a_974_n21642# A6 a_578_n21642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8414 GND A1 word360 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8415 word776 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8416 GND A3 word852 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8417 GND A8 word45 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8418 GND A0 word960 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8419 word333 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8420 word263 a_2376_n66# a_2162_n37546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8421 a_446_n34280# A8 a_182_n34280# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8422 a_1766_n16388# A3 a_1370_n16388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8423 a_974_n1194# A6 a_710_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8424 GND A1 word357 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8425 GND A8 word694 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8426 GND A0 word1016 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8427 GND A2 word425 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8428 GND A7 word606 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8429 GND A8 word764 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8430 word895 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8431 a_1766_n94062# A3 a_1370_n94062# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8432 GND A7 word547 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8433 a_2294_n119480# A1 a_2030_n119480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8434 a_974_n626# A6 a_710_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8435 a_578_n20222# a_528_n66# a_446_n20222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8436 a_182_n19512# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8437 GND A5 word13 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8438 GND A7 word64 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8439 GND A2 word323 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8440 word825 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8441 a_578_n58704# a_528_n66# a_314_n58704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8442 GND A2 word264 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8443 GND A6 word446 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8444 a_578_n139076# a_528_n66# a_314_n139076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8445 a_446_n89092# A8 a_50_n89092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8446 a_446_n9572# A8 a_182_n9572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8447 word540 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8448 word529 a_2376_n66# a_2294_n75318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8449 word950 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8450 a_50_n115930# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8451 a_50_n124308# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8452 a_974_n36552# A6 a_710_n36552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8453 GND A0 word448 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8454 GND A1 word465 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8455 GND A7 word325 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8456 word11 a_2376_n66# a_2162_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8457 a_2162_n5596# a_2112_n66# a_1898_n5596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8458 word957 a_2376_n66# a_2294_n136094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8459 word746 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8460 a_182_n10424# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8461 a_1370_n75886# a_1320_n66# a_1238_n75886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8462 a_1370_n84264# a_1320_n66# a_1238_n84264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8463 GND A6 word165 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8464 a_842_n67934# a_792_n66# a_578_n67934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8465 word167 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8466 word1012 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8467 GND A8 word528 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8468 GND A0 word346 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8469 word727 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8470 word959 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8471 a_1898_n31724# a_1848_n66# a_1634_n31724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8472 word377 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8473 word436 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8474 a_182_n48906# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8475 a_50_n123882# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8476 GND A1 word521 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8477 GND A2 word530 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8478 a_1502_n142058# A4 a_1106_n142058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8479 GND A5 word923 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8480 a_1106_n43084# a_1056_n66# a_974_n43084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8481 GND A2 word729 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8482 GND A6 word653 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8483 a_1502_n133680# A4 a_1106_n133680# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8484 a_578_n35132# a_528_n66# a_446_n35132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8485 a_578_n26754# a_528_n66# a_446_n26754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8486 GND A4 word160 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8487 a_842_n106842# a_792_n66# a_578_n106842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8488 a_842_n36410# a_792_n66# a_578_n36410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8489 word431 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8490 a_974_n74324# A6 a_710_n74324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8491 GND A8 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8492 GND A6 word551 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8493 a_2294_n2472# A1 a_2030_n2472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8494 word155 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8495 word245 a_2376_n66# a_2294_n34990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8496 GND A7 word100 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8497 GND A0 word282 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8498 word953 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8499 a_1502_n119196# A4 a_1238_n119196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8500 GND A1 word240 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8501 a_314_n46918# a_264_n66# a_182_n46918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8502 a_50_n139218# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8503 GND A0 word612 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8504 GND A0 word840 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8505 a_1766_n69070# A3 a_1502_n69070# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8506 word934 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8507 a_842_n35984# a_792_n66# a_578_n35984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8508 GND A7 word588 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8509 word846 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8510 word211 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8511 GND A4 word546 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8512 a_1370_n99174# a_1320_n66# a_1106_n99174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8513 a_182_n16956# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8514 a_182_n25334# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8515 word152 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8516 GND A6 word270 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8517 a_1106_n72478# a_1056_n66# a_842_n72478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8518 a_578_n64526# a_528_n66# a_314_n64526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8519 a_1898_n46634# a_1848_n66# a_1766_n46634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8520 GND A6 word428 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8521 word541 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8522 a_842_n144614# a_792_n66# a_578_n144614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8523 a_50_n86820# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8524 a_50_n138792# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8525 word37 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8526 a_2294_n9430# A1 a_2030_n9430# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8527 GND A5 word969 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8528 GND A2 word834 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8529 a_50_n130130# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8530 a_974_n42374# A6 a_710_n42374# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8531 word543 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8532 word762 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8533 GND A4 word324 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8534 GND A4 word265 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8535 word355 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8536 a_842_n82134# a_792_n66# a_710_n82134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8537 a_1370_n90086# a_1320_n66# a_1106_n90086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8538 a_50_n94772# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8539 word409 a_2376_n66# a_2294_n58278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8540 word477 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8541 a_50_n107268# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8542 word1000 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8543 a_182_n63106# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8544 GND A0 word328 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8545 GND A1 word345 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8546 a_182_n54728# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8547 a_1502_n36836# A4 a_1238_n36836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8548 GND A4 word321 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8549 a_578_n93920# a_528_n66# a_446_n93920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8550 word951 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8551 word984 A0 a_2294_n139928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8552 word892 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8553 a_842_n121042# a_792_n66# a_710_n121042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8554 a_578_n32576# a_528_n66# a_446_n32576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8555 a_1898_n14684# a_1848_n66# a_1766_n14684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8556 word316 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8557 word255 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8558 a_974_n80146# A6 a_710_n80146# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8559 a_1106_n87388# a_1056_n66# a_842_n87388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8560 a_182_n5028# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8561 GND A6 word533 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8562 word994 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8563 a_314_n61118# a_264_n66# a_182_n61118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8564 word935 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8565 a_314_n52740# a_264_n66# a_182_n52740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8566 GND A4 word99 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8567 word675 a_2376_n66# a_2162_n96050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8568 a_50_n145040# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8569 a_974_n116924# A6 a_710_n116924# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8570 a_842_n50184# a_792_n66# a_710_n50184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8571 word311 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8572 a_1634_n47202# a_1584_n66# a_1502_n47202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8573 a_974_n57284# A6 a_578_n57284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8574 GND A0 word594 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8575 word252 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8576 a_1502_n74608# A4 a_1238_n74608# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8577 word920 A0 a_2294_n130840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8578 a_314_n38256# a_264_n66# a_182_n38256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8579 GND A4 word587 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8580 word460 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8581 a_182_n22778# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8582 a_182_n31156# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8583 a_314_n60692# a_264_n66# a_182_n60692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8584 a_842_n88666# a_792_n66# a_710_n88666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8585 word151 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8586 a_578_n70348# a_528_n66# a_314_n70348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8587 word814 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8588 a_182_n69638# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8589 a_578_n61970# a_528_n66# a_314_n61970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8590 word726 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8591 word818 A0 a_2162_n116356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8592 word212 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8593 GND A2 word875 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8594 word584 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8595 word803 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8596 word744 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8597 word293 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8598 GND A4 word365 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8599 word525 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8600 a_50_n78158# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8601 a_1898_n29594# a_1848_n66# a_1634_n29594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8602 a_1238_n37404# A5 a_974_n37404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8603 a_974_n95056# A6 a_578_n95056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8604 word518 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8605 GND A6 word697 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8606 a_50_n113090# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8607 a_2162_n20932# a_2112_n66# a_2030_n20932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8608 word191 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8609 a_314_n67650# a_264_n66# a_182_n67650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8610 a_1634_n15252# a_1584_n66# a_1502_n15252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8611 a_1502_n51036# A4 a_1106_n51036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8612 a_1106_n134106# a_1056_n66# a_974_n134106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8613 a_182_n60550# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8614 GND A4 word204 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8615 a_1502_n42658# A4 a_1106_n42658# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8616 a_314_n122320# a_264_n66# a_50_n122320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8617 a_1106_n125728# a_1056_n66# a_842_n125728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8618 a_1634_n117918# a_1584_n66# a_1370_n117918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8619 a_1898_n105422# a_1848_n66# a_1766_n105422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8620 a_1502_n2330# A4 a_1238_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8621 a_842_n65094# a_792_n66# a_578_n65094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8622 word147 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8623 a_1898_n81850# a_1848_n66# a_1634_n81850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8624 GND A5 word143 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8625 word933 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8626 a_182_n46066# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8627 a_182_n37688# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8628 GND A2 word56 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8629 a_1502_n19796# A4 a_1238_n19796# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8630 a_1502_n28174# A4 a_1238_n28174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8631 word1010 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8632 a_3820_164# A3 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X8633 a_314_n130272# a_264_n66# a_50_n130272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8634 word418 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8635 word978 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8636 a_1898_n58988# a_1848_n66# a_1634_n58988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8637 a_314_n121894# a_264_n66# a_50_n121894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8638 word681 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8639 word628 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8640 GND A4 word140 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8641 GND A3 word532 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8642 word135 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8643 word908 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8644 a_1766_n134532# A3 a_1370_n134532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8645 a_974_n131124# A6 a_578_n131124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8646 word689 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8647 a_1634_n44646# a_1584_n66# a_1370_n44646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8648 word630 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8649 a_314_n44078# a_264_n66# a_182_n44078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8650 word98 A0 a_2162_n14116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8651 a_1898_n134816# a_1848_n66# a_1766_n134816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8652 a_1370_n3040# a_1320_n66# a_1238_n3040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8653 a_2162_n35842# a_2112_n66# a_2030_n35842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8654 word623 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8655 GND A3 word310 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8656 a_314_n137230# a_264_n66# a_50_n137230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8657 word586 A0 a_2162_n83412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8658 word564 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8659 a_1766_n103008# A3 a_1370_n103008# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8660 word684 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8661 word340 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8662 word800 A0 a_2294_n113800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8663 word463 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8664 word522 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8665 word844 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8666 word785 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8667 GND A7 word831 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8668 GND A7 word772 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8669 GND A3 word307 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8670 GND A9 word241 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8671 a_2294_n33854# A1 a_1898_n33854# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8672 word92 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8673 a_2294_n42232# A1 a_2030_n42232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8674 a_314_n145182# a_264_n66# a_50_n145182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8675 a_974_n92500# A6 a_578_n92500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8676 a_1766_n102582# A3 a_1370_n102582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8677 a_1634_n12696# a_1584_n66# a_1370_n12696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8678 word173 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8679 GND A8 word81 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8680 word991 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8681 word706 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8682 GND A1 word836 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8683 a_446_n104712# A8 a_50_n104712# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8684 a_1898_n111244# a_1848_n66# a_1634_n111244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8685 word234 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8686 a_710_n77732# A7 a_446_n77732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8687 GND A3 word85 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8688 word977 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8689 a_1106_n117066# a_1056_n66# a_974_n117066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8690 a_1106_n108688# a_1056_n66# a_842_n108688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8691 a_2030_n111528# A2 a_1766_n111528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8692 GND A5 word455 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8693 word400 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8694 word459 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8695 a_1634_n131692# a_1584_n66# a_1370_n131692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8696 word238 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8697 a_578_n91080# a_528_n66# a_446_n91080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8698 word669 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8699 word632 A0 a_2294_n89944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8700 GND A9 word448 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8701 word964 A0 a_2294_n137088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8702 a_1238_n11276# A5 a_842_n11276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8703 word627 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8704 a_1766_n109540# A3 a_1502_n109540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8705 a_710_n46208# A7 a_314_n46208# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8706 word358 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8707 a_1766_n131976# A3 a_1502_n131976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8708 a_710_n37830# A7 a_314_n37830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8709 a_2030_n19938# A2 a_1634_n19938# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8710 word439 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8711 word890 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8712 word755 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8713 a_1238_n58136# A5 a_974_n58136# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8714 word561 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8715 a_2162_n104428# a_2112_n66# a_1898_n104428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8716 word80 A0 a_2294_n11560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8717 a_1238_n49758# A5 a_842_n49758# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8718 GND A3 word471 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8719 word629 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8720 GND A9 word346 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8721 a_2162_n19228# a_2112_n66# a_1898_n19228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8722 a_2294_n57142# A1 a_2030_n57142# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8723 a_1634_n97328# a_1584_n66# a_1502_n97328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8724 a_1898_n140638# a_1848_n66# a_1634_n140638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8725 a_2162_n50042# a_2112_n66# a_1898_n50042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8726 word197 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8727 a_974_n114084# A6 a_710_n114084# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8728 word337 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8729 word410 A0 a_2162_n58420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8730 a_710_n45782# A7 a_314_n45782# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8731 a_4612_164# A6 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X8732 GND A8 word186 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8733 word568 A0 a_2294_n80856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8734 a_2162_n88524# a_2112_n66# a_1898_n88524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8735 a_1634_n138650# a_1584_n66# a_1502_n138650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8736 word752 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8737 a_1898_n126154# a_1848_n66# a_1766_n126154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8738 word563 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8739 a_1898_n117776# a_1848_n66# a_1634_n117776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8740 a_2030_n10850# A2 a_1634_n10850# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8741 word497 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8742 GND A7 word872 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8743 a_1238_n40670# A5 a_974_n40670# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8744 word466 A0 a_2162_n66372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8745 GND A7 word813 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8746 a_2030_n126438# A2 a_1634_n126438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8747 a_2162_n10140# a_2112_n66# a_1898_n10140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8748 a_2294_n17240# A1 a_2030_n17240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8749 GND A9 word282 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8750 GND A9 word223 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8751 word402 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8752 a_710_n14258# A7 a_446_n14258# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8753 word91 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8754 GND A5 word128 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8755 GND A3 word678 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8756 a_2294_n86536# A1 a_2030_n86536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8757 GND A1 word936 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8758 GND A3 word881 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8759 GND A1 word877 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8760 GND A9 word121 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8761 word881 a_2376_n66# a_2294_n125302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8762 GND A3 word822 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8763 a_2294_n25192# A1 a_2030_n25192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8764 a_1634_n65378# a_1584_n66# a_1502_n65378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8765 a_710_n83554# A7 a_446_n83554# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8766 a_2162_n119338# a_2112_n66# a_1898_n119338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8767 a_1238_n95482# A5 a_974_n95482# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8768 word1018 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8769 word786 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8770 a_1634_n106700# a_1584_n66# a_1502_n106700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8771 a_1370_n122604# a_1320_n66# a_1238_n122604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8772 a_1634_n115078# a_1584_n66# a_1502_n115078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8773 a_974_n5312# A6 a_710_n5312# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8774 word500 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8775 GND A9 word62 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8776 word11 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8777 word114 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8778 a_1502_n78300# A4 a_1106_n78300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8779 a_1106_n23914# a_1056_n66# a_974_n23914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8780 a_710_n52030# A7 a_314_n52030# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8781 GND A8 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8782 a_1766_n89802# A3 a_1370_n89802# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8783 GND A5 word394 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8784 word298 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8785 GND A5 word335 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8786 a_2162_n110250# a_2112_n66# a_1898_n110250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8787 a_1238_n55580# A5 a_974_n55580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8788 word1012 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8789 GND A9 word387 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8790 a_2162_n25050# a_2112_n66# a_1898_n25050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8791 GND A9 word328 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8792 GND A4 word941 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8793 word979 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8794 word137 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8795 word319 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8796 GND A8 word227 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8797 a_2162_n94346# a_2112_n66# a_1898_n94346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8798 word717 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8799 GND A7 word512 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8800 GND A8 word729 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8801 word852 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8802 a_2162_n9714# a_2112_n66# a_2030_n9714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8803 a_1766_n80714# A3 a_1370_n80714# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8804 a_1238_n128852# A5 a_974_n128852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8805 a_1898_n123598# a_1848_n66# a_1766_n123598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8806 a_2294_n114510# A1 a_1898_n114510# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8807 word380 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8808 GND A7 word29 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8809 word891 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8810 GND A7 word854 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8811 a_2030_n132260# A2 a_1766_n132260# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8812 a_578_n134106# a_528_n66# a_314_n134106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8813 word976 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8814 a_446_n4602# A8 a_182_n4602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8815 a_446_n84122# A8 a_50_n84122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8816 word857 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8817 a_446_n75744# A8 a_50_n75744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8818 a_1766_n57852# A3 a_1370_n57852# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8819 word505 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8820 word915 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8821 a_2294_n122462# A1 a_1898_n122462# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8822 GND A1 word760 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8823 word73 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8824 a_2294_n92358# A1 a_2030_n92358# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8825 GND A7 word26 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8826 a_2030_n49048# A2 a_1634_n49048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8827 a_2030_n109398# A2 a_1766_n109398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8828 word787 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8829 word846 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8830 word585 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8831 GND A4 word716 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8832 word863 a_2376_n66# a_2162_n122746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8833 a_710_n80998# A7 a_446_n80998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8834 a_1370_n70916# a_1320_n66# a_1106_n70916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8835 GND A5 word657 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8836 word754 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8837 word924 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8838 GND A1 word816 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8839 a_2162_n62396# a_2112_n66# a_1898_n62396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8840 a_2294_n69496# A1 a_2030_n69496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8841 GND A7 word287 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8842 GND A1 word757 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8843 a_974_n2756# A6 a_710_n2756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8844 word761 a_2376_n66# a_2294_n108262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8845 GND A9 word44 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8846 word965 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8847 GND A7 word617 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8848 word763 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8849 a_578_n102156# a_528_n66# a_446_n102156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8850 word650 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8851 a_1766_n95624# A3 a_1502_n95624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8852 GND A5 word24 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8853 word181 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8854 word485 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8855 word921 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8856 GND A2 word393 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8857 a_1502_n114226# A4 a_1106_n114226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8858 GND A5 word727 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8859 a_1106_n15252# a_1056_n66# a_842_n15252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8860 a_1502_n105848# A4 a_1106_n105848# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8861 word1021 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8862 GND A9 word369 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8863 a_446_n99032# A8 a_50_n99032# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8864 a_1370_n16530# a_1320_n66# a_1106_n16530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8865 word1020 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8866 word951 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8867 GND A0 word86 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8868 word892 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8869 a_446_n12270# A8 a_182_n12270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8870 a_1370_n94204# a_1320_n66# a_1238_n94204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8871 a_710_n110392# A7 a_314_n110392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8872 a_1370_n85826# a_1320_n66# a_1238_n85826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8873 GND A8 word598 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8874 GND A8 word539 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8875 word666 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8876 a_1370_n143336# a_1320_n66# a_1106_n143336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8877 word970 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8878 GND A8 word107 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8879 a_1370_n134958# a_1320_n66# a_1106_n134958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8880 a_578_n131550# a_528_n66# a_314_n131550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8881 a_50_n133822# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8882 word29 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8883 GND A1 word532 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8884 a_446_n81566# A8 a_50_n81566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8885 GND A2 word168 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8886 a_1106_n44646# a_1056_n66# a_974_n44646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8887 a_1106_n53024# a_1056_n66# a_842_n53024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8888 a_1238_n103150# A5 a_842_n103150# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8889 GND A6 word291 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8890 a_578_n108688# a_528_n66# a_446_n108688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8891 word444 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8892 GND A5 word832 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8893 word26 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8894 word315 a_2376_n66# a_2162_n44930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8895 a_1502_n129136# A4 a_1238_n129136# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8896 GND A5 word773 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8897 a_710_n117350# A7 a_314_n117350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8898 GND A2 word656 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8899 GND A3 word802 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8900 a_1766_n32150# A3 a_1502_n32150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8901 GND A0 word910 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8902 a_842_n54302# a_792_n66# a_710_n54302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8903 a_1370_n53876# a_1320_n66# a_1106_n53876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8904 a_1370_n62254# a_1320_n66# a_1106_n62254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8905 a_842_n45924# a_792_n66# a_710_n45924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8906 word745 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8907 a_446_n27180# A8 a_182_n27180# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8908 GND A0 word132 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8909 word222 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8910 word281 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8911 word371 a_2376_n66# a_2162_n52882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8912 a_50_n101872# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8913 a_1370_n39392# a_1320_n66# a_1238_n39392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8914 GND A0 word966 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8915 GND A4 word865 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8916 word843 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8917 a_1502_n120048# A4 a_1238_n120048# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8918 GND A5 word709 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8919 GND A1 word696 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8920 word701 a_2376_n66# a_2294_n99742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8921 GND A7 word556 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8922 a_446_n96476# A8 a_50_n96476# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8923 word219 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8924 word149 a_2376_n66# a_2294_n21358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8925 a_974_n43936# A6 a_710_n43936# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8926 a_1106_n59556# a_1056_n66# a_974_n59556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8927 GND A6 word396 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8928 GND A3 word1009 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8929 word992 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8930 word933 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8931 word1009 a_2376_n66# a_2294_n143478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8932 a_1238_n140496# A5 a_842_n140496# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8933 GND A1 word85 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8934 a_710_n6874# A7 a_446_n6874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8935 word479 a_2376_n66# a_2162_n68218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8936 word490 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8937 GND A8 word580 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8938 a_50_n117208# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8939 GND A7 word275 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8940 a_50_n108830# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8941 GND A0 word398 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8942 word637 a_2376_n66# a_2294_n90654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8943 a_1370_n140780# a_1320_n66# a_1238_n140780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8944 word779 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8945 a_842_n13974# a_792_n66# a_710_n13974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8946 GND A1 word573 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8947 GND A4 word391 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8948 a_1370_n77164# a_1320_n66# a_1238_n77164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8949 a_842_n69212# a_792_n66# a_578_n69212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8950 a_1106_n50468# a_1056_n66# a_842_n50468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8951 word909 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8952 a_1370_n126296# a_1320_n66# a_1106_n126296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8953 a_1898_n24624# a_1848_n66# a_1634_n24624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8954 a_1898_n33002# a_1848_n66# a_1766_n33002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8955 a_842_n122604# a_792_n66# a_710_n122604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8956 a_50_n116782# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8957 a_974_n81708# A6 a_710_n81708# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8958 a_1106_n97328# a_1056_n66# a_974_n97328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8959 GND A2 word480 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8960 a_1106_n88950# a_1056_n66# a_842_n88950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8961 GND A6 word662 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8962 a_974_n20364# A6 a_578_n20364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8963 word1005 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8964 a_578_n19654# a_528_n66# a_446_n19654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8965 a_578_n28032# a_528_n66# a_446_n28032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8966 GND A6 word171 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8967 GND A4 word110 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8968 a_842_n29310# a_792_n66# a_578_n29310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8969 word381 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8970 a_842_n51746# a_792_n66# a_710_n51746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8971 a_974_n58846# A6 a_578_n58846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8972 word845 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8973 word195 a_2376_n66# a_2162_n27890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8974 GND A0 word232 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8975 a_182_n32718# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8976 a_314_n39818# a_264_n66# a_182_n39818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8977 a_1502_n23204# A4 a_1106_n23204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8978 a_314_n70632# a_264_n66# a_182_n70632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8979 a_1502_n14826# A4 a_1106_n14826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8980 GND A8 word685 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8981 GND A4 word166 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8982 word1019 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8983 word943 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8984 a_842_n28884# a_792_n66# a_578_n28884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8985 a_578_n71910# a_528_n66# a_314_n71910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8986 word593 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8987 GND A7 word538 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8988 word796 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8989 a_182_n18234# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8990 GND A6 word437 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8991 a_842_n137514# a_792_n66# a_578_n137514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8992 a_578_n57426# a_528_n66# a_314_n57426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8993 a_1898_n39534# a_1848_n66# a_1766_n39534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8994 a_446_n8294# A8 a_182_n8294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8995 a_50_n79720# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8996 GND A4 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X8997 GND A3 word336 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X8998 a_974_n96618# A6 a_578_n96618# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X8999 GND A5 word978 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9000 a_50_n123030# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9001 a_974_n26896# A6 a_578_n26896# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9002 word156 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9003 GND A2 word1001 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9004 GND A6 word276 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9005 word651 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9006 word305 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9007 a_50_n87672# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9008 word486 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9009 word217 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9010 a_842_n66656# a_792_n66# a_578_n66656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9011 word158 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9012 word718 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9013 a_1898_n30446# a_1848_n66# a_1766_n30446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9014 GND A0 word278 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9015 a_182_n47628# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9016 a_182_n56006# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9017 GND A2 word67 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9018 a_1502_n38114# A4 a_1238_n38114# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9019 word368 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9020 a_314_n140212# a_264_n66# a_50_n140212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9021 GND A4 word271 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9022 a_314_n131834# a_264_n66# a_50_n131834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9023 a_1898_n77306# a_1848_n66# a_1634_n77306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9024 GND A2 word720 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9025 GND A6 word644 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9026 word646 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9027 word361 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9028 a_1898_n68928# a_1848_n66# a_1766_n68928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9029 word698 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9030 word901 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9031 a_578_n25476# a_528_n66# a_446_n25476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9032 a_842_n105564# a_792_n66# a_578_n105564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9033 word13 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9034 word205 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9035 word422 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9036 a_974_n73046# A6 a_710_n73046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9037 word295 a_2376_n66# a_2162_n42090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9038 GND A6 word542 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9039 word944 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9040 a_314_n45640# a_264_n66# a_182_n45640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9041 a_314_n54018# a_264_n66# a_182_n54018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9042 GND A0 word214 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9043 a_578_n94772# a_528_n66# a_446_n94772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9044 word885 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9045 GND A2 word776 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9046 word693 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9047 word424 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9048 a_974_n118202# A6 a_710_n118202# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9049 a_974_n109824# A6 a_710_n109824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9050 word261 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9051 GND A0 word544 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9052 word634 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9053 a_1766_n5596# A3 a_1502_n5596# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9054 word575 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9055 word410 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9056 word870 A0 a_2162_n123740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9057 a_182_n24056# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9058 a_182_n15678# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9059 a_314_n53592# a_264_n66# a_182_n53592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9060 word855 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9061 a_1106_n71200# a_1056_n66# a_842_n71200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9062 a_842_n143336# a_792_n66# a_578_n143336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9063 word823 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9064 a_578_n54870# a_528_n66# a_314_n54870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9065 a_578_n63248# a_528_n66# a_314_n63248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9066 a_1898_n45356# a_1848_n66# a_1634_n45356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9067 word473 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9068 word768 A0 a_2294_n109256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9069 word414 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9070 GND A3 word436 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9071 word926 A0 a_2162_n131692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9072 word103 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9073 word753 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9074 word466 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9075 word407 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9076 GND A2 word825 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9077 a_1766_n112522# A3 a_1370_n112522# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9078 a_710_n40812# A7 a_314_n40812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9079 a_1634_n22636# a_1584_n66# a_1370_n22636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9080 a_1634_n31014# a_1584_n66# a_1370_n31014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9081 word243 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9082 a_974_n41096# A6 a_710_n41096# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9083 word534 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9084 word59 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9085 a_50_n93494# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9086 word468 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9087 a_974_n79578# A6 a_710_n79578# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9088 word527 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9089 a_842_n72478# a_792_n66# a_578_n72478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9090 a_182_n53450# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9091 a_314_n115220# a_264_n66# a_50_n115220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9092 word704 A0 a_2294_n100168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9093 a_1106_n127006# a_1056_n66# a_842_n127006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9094 word367 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9095 word470 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9096 GND A5 word93 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9097 a_1898_n74750# a_1848_n66# a_1634_n74750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9098 a_578_n31298# a_528_n66# a_446_n31298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9099 a_1238_n21216# A5 a_974_n21216# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9100 word301 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9101 GND A3 word643 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9102 a_1238_n12838# A5 a_842_n12838# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9103 a_1766_n141916# A3 a_1502_n141916# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9104 GND A3 word211 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9105 word960 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9106 GND A9 word86 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9107 a_2294_n20222# A1 a_1898_n20222# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9108 word206 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9109 a_1634_n60408# a_1584_n66# a_1502_n60408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9110 a_314_n114794# a_264_n66# a_50_n114794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9111 a_314_n123172# a_264_n66# a_50_n123172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9112 word631 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9113 word77 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9114 a_578_n69780# a_528_n66# a_314_n69780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9115 GND A5 word581 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9116 GND A3 word64 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9117 GND A3 word482 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9118 a_2162_n51604# a_2112_n66# a_2030_n51604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9119 a_2294_n58704# A1 a_1898_n58704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9120 a_1634_n101730# a_1584_n66# a_1502_n101730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9121 a_1766_n127432# A3 a_1502_n127432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9122 word302 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9123 word208 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9124 a_974_n115646# A6 a_710_n115646# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9125 word1016 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9126 a_1502_n73330# A4 a_1238_n73330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9127 word881 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9128 word54 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9129 GND A4 word519 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9130 word574 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9131 GND A4 word578 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9132 a_182_n21500# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9133 a_842_n87388# a_792_n66# a_710_n87388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9134 word142 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9135 word245 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9136 word83 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9137 GND A3 word260 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9138 a_1898_n42800# a_1848_n66# a_1634_n42800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9139 a_1898_n51178# a_1848_n66# a_1766_n51178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9140 word567 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9141 a_842_n140780# a_792_n66# a_578_n140780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9142 a_182_n68360# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9143 word536 A0 a_2294_n76312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9144 word750 A0 a_2162_n106700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9145 GND A9 word293 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9146 a_1898_n89660# a_1848_n66# a_1766_n89660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9147 word507 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9148 a_710_n15820# A7 a_446_n15820# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9149 GND A5 word139 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9150 GND A5 word198 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9151 word735 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9152 a_842_n126296# a_792_n66# a_710_n126296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9153 a_1238_n27748# A5 a_842_n27748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9154 word474 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9155 GND A9 word191 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9156 GND A3 word257 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9157 a_314_n138082# a_264_n66# a_50_n138082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9158 word509 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9159 GND A9 word132 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9160 a_2030_n75602# A2 a_1766_n75602# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9161 word123 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9162 a_1502_n41380# A4 a_1106_n41380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9163 word941 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9164 a_1634_n125018# a_1584_n66# a_1502_n125018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9165 a_1106_n124450# a_1056_n66# a_842_n124450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9166 a_2162_n66514# a_2112_n66# a_2030_n66514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9167 a_1898_n104144# a_1848_n66# a_1634_n104144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9168 GND A0 word690 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9169 word184 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9170 a_1502_n88240# A4 a_1106_n88240# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9171 GND A6 word805 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9172 GND A5 word75 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9173 word125 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9174 a_1634_n74892# a_1584_n66# a_1502_n74892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9175 word611 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9176 GND A4 word683 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9177 GND A3 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9178 word679 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9179 a_2162_n128852# a_2112_n66# a_2030_n128852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9180 word252 A0 a_2294_n35984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9181 word409 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9182 word247 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9183 GND A5 word405 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9184 word672 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9185 a_1634_n124592# a_1584_n66# a_1502_n124592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9186 a_1238_n65520# A5 a_842_n65520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9187 a_1502_n96192# A4 a_1106_n96192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9188 GND A9 word398 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9189 a_2294_n64526# A1 a_1898_n64526# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9190 GND A1 word781 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9191 a_710_n39108# A7 a_314_n39108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9192 word249 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9193 word840 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9194 a_2030_n43652# A2 a_1766_n43652# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9195 word389 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9196 GND A5 word461 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9197 word863 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9198 a_1238_n73472# A5 a_974_n73472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9199 a_2162_n95908# a_2112_n66# a_2030_n95908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9200 word614 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9201 word716 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9202 a_2162_n34564# a_2112_n66# a_2030_n34564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9203 a_1766_n20932# A3 a_1370_n20932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9204 a_710_n38682# A7 a_314_n38682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9205 a_1502_n56290# A4 a_1238_n56290# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9206 word518 A0 a_2162_n73756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9207 word675 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9208 word761 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9209 word24 A0 a_2294_n3608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9210 GND A8 word136 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9211 word927 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9212 a_1898_n119054# a_1848_n66# a_1766_n119054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9213 GND A0 word14 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9214 word454 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9215 word506 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9216 GND A6 word910 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9217 a_446_n15962# A8 a_182_n15962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9218 word143 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9219 word447 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9220 a_1106_n6306# a_1056_n66# a_974_n6306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9221 word416 A0 a_2294_n59272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9222 a_2294_n93920# A1 a_1898_n93920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9223 GND A9 word232 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9224 a_1634_n81140# a_1584_n66# a_1370_n81140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9225 word655 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9226 GND A9 word173 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9227 a_2294_n32576# A1 a_1898_n32576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9228 a_710_n90938# A7 a_446_n90938# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9229 word765 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9230 a_1238_n19086# A5 a_974_n19086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9231 GND A3 word628 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9232 word705 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9233 GND A8 word72 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9234 GND A6 word907 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9235 a_1766_n139786# A3 a_1370_n139786# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9236 a_974_n136378# A6 a_578_n136378# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9237 GND A3 word772 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9238 a_446_n103434# A8 a_50_n103434# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9239 a_974_n128000# A6 a_578_n128000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9240 word831 a_2376_n66# a_2162_n118202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9241 word225 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9242 a_1634_n49900# a_1584_n66# a_1370_n49900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9243 a_710_n76454# A7 a_446_n76454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9244 a_1634_n58278# a_1584_n66# a_1370_n58278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9245 a_2030_n58562# A2 a_1634_n58562# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9246 word968 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9247 a_2162_n143052# a_2112_n66# a_1898_n143052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9248 a_2162_n134674# a_2112_n66# a_2030_n134674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9249 GND A2 word74 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9250 word352 A0 a_2294_n50184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9251 a_578_n103718# a_528_n66# a_446_n103718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9252 word555 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9253 word450 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9254 word991 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9255 GND A1 word336 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9256 a_2162_n49474# a_2112_n66# a_2030_n49474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9257 word682 A0 a_2162_n97044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9258 GND A3 word564 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9259 GND A9 word439 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9260 a_1106_n16814# a_1056_n66# a_842_n16814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9261 word559 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9262 a_2030_n18660# A2 a_1766_n18660# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9263 GND A5 word344 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9264 GND A3 word708 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9265 a_2294_n138934# A1 a_2030_n138934# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9266 a_1766_n130698# A3 a_1370_n130698# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9267 GND A1 word61 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9268 word248 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9269 a_1238_n48480# A5 a_842_n48480# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9270 word552 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9271 word620 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9272 word962 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9273 GND A9 word337 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9274 GND A9 word278 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9275 a_446_n22210# A8 a_182_n22210# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9276 a_710_n120332# A7 a_314_n120332# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9277 a_2162_n40386# a_2112_n66# a_2030_n40386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9278 a_2294_n47486# A1 a_1898_n47486# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9279 a_2030_n87956# A2 a_1634_n87956# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9280 a_710_n111954# A7 a_314_n111954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9281 a_182_n768# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9282 word269 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9283 GND A8 word16 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9284 a_1370_n34422# a_1320_n66# a_1106_n34422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9285 GND A8 word177 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9286 GND A8 word118 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9287 a_2162_n78868# a_2112_n66# a_2030_n78868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9288 word495 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9289 a_1766_n73614# A3 a_1502_n73614# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9290 a_446_n91506# A8 a_50_n91506# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9291 a_446_n21784# A8 a_182_n21784# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9292 a_446_n30162# A8 a_182_n30162# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9293 GND A6 word47 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9294 GND A7 word804 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9295 a_3028_164# A0 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X9296 GND A2 word179 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9297 a_2030_n125160# A2 a_1766_n125160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9298 a_446_n77022# A8 a_50_n77022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9299 GND A9 word214 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9300 word807 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9301 a_710_n1904# A7 a_446_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9302 a_2294_n106984# A1 a_2030_n106984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9303 GND A5 word843 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9304 GND A8 word65 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9305 a_2294_n76880# A1 a_1898_n76880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9306 GND A2 word667 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9307 word796 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9308 GND A1 word868 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9309 a_1238_n121042# A5 a_842_n121042# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9310 a_446_n100878# A8 a_50_n100878# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9311 word535 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9312 word813 a_2376_n66# a_2294_n115646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9313 a_1238_n112664# A5 a_974_n112664# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9314 a_710_n73898# A7 a_446_n73898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9315 a_710_n82276# A7 a_446_n82276# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9316 a_2162_n118060# a_2112_n66# a_1898_n118060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9317 GND A5 word607 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9318 word1009 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9319 word511 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9320 GND A0 word706 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9321 word874 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9322 a_1370_n121326# a_1320_n66# a_1238_n121326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9323 word815 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9324 a_1766_n19228# A3 a_1502_n19228# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9325 word441 a_2376_n66# a_2294_n62822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9326 GND A7 word296 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9327 a_1370_n112948# a_1320_n66# a_1238_n112948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9328 a_974_n4034# A6 a_710_n4034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9329 a_50_n111812# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9330 GND A1 word377 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9331 GND A1 word436 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9332 a_710_n126864# A7 a_314_n126864# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9333 a_1766_n41664# A3 a_1502_n41664# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9334 a_1370_n49332# a_1320_n66# a_1238_n49332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9335 GND A5 word779 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9336 word664 A0 a_2294_n94488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9337 word1003 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9338 GND A9 word319 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9339 word971 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9340 a_1766_n10140# A3 a_1502_n10140# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9341 GND A2 word442 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9342 GND A4 word932 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9343 a_2030_n93778# A2 a_1766_n93778# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9344 a_1370_n31866# a_1320_n66# a_1238_n31866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9345 a_1370_n40244# a_1320_n66# a_1238_n40244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9346 GND A8 word218 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9347 GND A7 word562 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9348 GND A8 word720 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9349 word31 a_2376_n66# a_2162_n4602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9350 a_2162_n8436# a_2112_n66# a_2030_n8436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9351 GND A8 word159 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9352 a_2162_n84690# a_2112_n66# a_2030_n84690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9353 a_2162_n93068# a_2112_n66# a_1898_n93068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9354 word842 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9355 word901 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9356 GND A1 word973 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9357 a_1238_n127574# A5 a_974_n127574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9358 GND A4 word771 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9359 GND A7 word20 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9360 GND A7 word71 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9361 GND A8 word548 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9362 GND A1 word152 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9363 a_1106_n60408# a_1056_n66# a_974_n60408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9364 word616 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9365 GND A7 word845 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9366 word882 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9367 a_1370_n17382# a_1320_n66# a_1106_n17382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9368 GND A4 word710 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9369 a_1370_n136236# a_1320_n66# a_1106_n136236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9370 a_2162_n484# a_2112_n66# a_2030_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9371 a_50_n126722# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9372 GND A7 word342 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9373 GND A1 word541 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9374 GND A0 word752 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9375 a_446_n3324# A8 a_182_n3324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9376 a_446_n74466# A8 a_50_n74466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9377 a_2294_n121184# A1 a_1898_n121184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9378 a_1502_n136520# A4 a_1238_n136520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9379 a_974_n21926# A6 a_578_n21926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9380 a_2294_n91080# A1 a_2030_n91080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9381 GND A3 word854 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9382 word778 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9383 word394 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9384 GND A4 word707 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9385 a_50_n82702# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9386 word335 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9387 a_2294_n5312# A1 a_1898_n5312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9388 GND A7 word120 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9389 word265 a_2376_n66# a_2294_n37830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9390 GND A1 word260 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9391 GND A2 word547 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9392 GND A9 word35 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9393 a_3820_164# A3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X9394 a_974_n1478# A6 a_710_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9395 GND A4 word236 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9396 a_842_n47202# a_792_n66# a_710_n47202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9397 GND A7 word608 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9398 GND A0 word1018 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9399 a_1766_n9714# A3 a_1502_n9714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9400 a_1766_n94346# A3 a_1370_n94346# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9401 a_1370_n104286# a_1320_n66# a_1238_n104286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9402 a_974_n910# A6 a_710_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9403 a_578_n20506# a_528_n66# a_446_n20506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9404 word321 a_2376_n66# a_2294_n45782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9405 GND A5 word15 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9406 GND A1 word316 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9407 GND A1 word257 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9408 GND A5 word718 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9409 a_578_n139360# a_528_n66# a_314_n139360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9410 word50 A0 a_2162_n7300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9411 a_446_n9856# A8 a_182_n9856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9412 a_446_n89376# A8 a_50_n89376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9413 a_2294_n136094# A1 a_1898_n136094# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9414 word169 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9415 a_974_n45214# A6 a_710_n45214# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9416 word99 a_2376_n66# a_2162_n14258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9417 word167 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9418 a_974_n36836# A6 a_710_n36836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9419 word883 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9420 GND A3 word900 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9421 word959 a_2376_n66# a_2162_n136378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9422 word748 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9423 a_182_n10708# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9424 a_710_n8152# A7 a_446_n8152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9425 a_50_n97612# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9426 a_1370_n84548# a_1320_n66# a_1238_n84548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9427 word1020 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9428 GND A8 word530 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9429 word923 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9430 GND A0 word348 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9431 word587 a_2376_n66# a_2162_n83554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9432 GND A0 word852 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9433 a_842_n15252# a_792_n66# a_710_n15252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9434 a_50_n132544# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9435 GND A7 word383 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9436 word20 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9437 a_446_n80288# A8 a_50_n80288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9438 a_1766_n62396# A3 a_1370_n62396# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9439 word431 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9440 GND A5 word925 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9441 a_578_n35416# a_528_n66# a_446_n35416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9442 a_1106_n34990# a_1056_n66# a_842_n34990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9443 a_1106_n43368# a_1056_n66# a_974_n43368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9444 GND A6 word282 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9445 word277 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9446 a_50_n109682# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9447 word24 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9448 GND A3 word181 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9449 word365 a_2376_n66# a_2294_n52030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9450 a_974_n74608# A6 a_710_n74608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9451 a_314_n118912# a_264_n66# a_50_n118912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9452 a_50_n101020# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9453 GND A6 word553 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9454 a_1502_n119480# A4 a_1238_n119480# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9455 a_1634_n1336# a_1584_n66# a_1502_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9456 GND A0 word284 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9457 word955 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9458 GND A2 word787 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9459 a_842_n53024# a_792_n66# a_710_n53024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9460 a_1370_n52598# a_1320_n66# a_1106_n52598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9461 GND A7 word590 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9462 word795 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9463 a_710_n200# A7 a_446_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9464 GND A0 word182 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9465 a_1766_n91790# A3 a_1502_n91790# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9466 a_182_n7442# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9467 a_182_n25618# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9468 a_50_n100594# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9469 word213 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9470 a_1370_n99458# a_1320_n66# a_1106_n99458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9471 word1011 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9472 a_314_n63532# a_264_n66# a_182_n63532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9473 a_1106_n81140# a_1056_n66# a_974_n81140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9474 a_578_n64810# a_528_n66# a_314_n64810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9475 word834 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9476 word543 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9477 word39 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9478 a_446_n95198# A8 a_50_n95198# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9479 GND A1 word628 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9480 word996 A0 a_2294_n141632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9481 word477 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9482 a_974_n42658# A6 a_710_n42658# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9483 GND A6 word387 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9484 a_578_n72762# a_528_n66# a_314_n72762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9485 a_1370_n90370# a_1320_n66# a_1106_n90370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9486 a_710_n5596# A7 a_446_n5596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9487 a_842_n82418# a_792_n66# a_710_n82418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9488 a_842_n12696# a_792_n66# a_710_n12696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9489 a_974_n19796# A6 a_578_n19796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9490 word569 a_2376_n66# a_2294_n80998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9491 word774 A0 a_2162_n110108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9492 GND A1 word564 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9493 word601 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9494 a_842_n121326# a_792_n66# a_710_n121326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9495 a_578_n32860# a_528_n66# a_446_n32860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9496 word318 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9497 a_842_n81992# a_792_n66# a_710_n81992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9498 a_182_n62964# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9499 a_182_n71342# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9500 a_974_n80430# A6 a_710_n80430# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9501 a_314_n124734# a_264_n66# a_50_n124734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9502 a_314_n133112# a_264_n66# a_50_n133112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9503 a_1106_n96050# a_1056_n66# a_974_n96050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9504 word311 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9505 a_578_n18376# a_528_n66# a_446_n18376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9506 a_1502_n4744# A4 a_1106_n4744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9507 a_842_n50468# a_792_n66# a_710_n50468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9508 a_974_n57568# A6 a_578_n57568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9509 word372 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9510 word894 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9511 GND A0 word164 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9512 GND A4 word648 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9513 a_182_n4886# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9514 a_182_n31440# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9515 a_314_n38540# a_264_n66# a_182_n38540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9516 GND A4 word589 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9517 a_314_n60976# a_264_n66# a_182_n60976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9518 a_842_n88950# a_792_n66# a_710_n88950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9519 a_1898_n61118# a_1848_n66# a_1634_n61118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9520 word875 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9521 word57 a_2376_n66# a_2294_n8294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9522 GND A1 word669 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9523 word820 A0 a_2294_n116640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9524 a_50_n144898# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9525 GND A4 word487 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9526 a_1502_n91222# A4 a_1238_n91222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9527 GND A0 word652 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9528 a_2030_n2898# A2 a_1766_n2898# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9529 word53 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9530 a_1502_n82844# A4 a_1238_n82844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9531 a_314_n46492# a_264_n66# a_182_n46492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9532 word805 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9533 a_578_n56148# a_528_n66# a_314_n56148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9534 a_1898_n38256# a_1848_n66# a_1634_n38256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9535 GND A3 word386 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9536 GND A3 word327 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9537 a_974_n95340# A6 a_578_n95340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9538 word876 A0 a_2294_n124592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9539 word112 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9540 a_1502_n59982# A4 a_1106_n59982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9541 a_314_n139644# a_264_n66# a_50_n139644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9542 a_1766_n105422# A3 a_1502_n105422# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9543 word416 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9544 GND A6 word699 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9545 GND A0 word430 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9546 word701 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9547 GND A2 word992 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9548 a_1634_n15536# a_1584_n66# a_1502_n15536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9549 word193 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9550 a_1502_n51320# A4 a_1106_n51320# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9551 word861 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9552 word583 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9553 word642 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9554 GND A4 word364 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9555 GND A4 word423 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9556 a_1898_n105706# a_1848_n66# a_1766_n105706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9557 a_50_n86394# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9558 a_842_n65378# a_792_n66# a_578_n65378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9559 word149 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9560 word681 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9561 word935 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9562 a_182_n46350# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9563 GND A2 word58 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9564 a_1502_n28458# A4 a_1238_n28458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9565 word322 A0 a_2162_n45924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9566 word479 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9567 a_1502_n50894# A4 a_1106_n50894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9568 a_314_n130556# a_264_n66# a_50_n130556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9569 word420 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9570 a_1106_n142342# a_1056_n66# a_842_n142342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9571 a_1106_n133964# a_1056_n66# a_974_n133964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9572 word258 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9573 a_1898_n76028# a_1848_n66# a_1766_n76028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9574 word689 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9575 word352 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9576 GND A3 word593 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9577 word630 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9578 a_578_n24198# a_528_n66# a_446_n24198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9579 word251 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9580 a_842_n104286# a_792_n66# a_578_n104286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9581 a_1502_n97754# A4 a_1106_n97754# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9582 GND A6 word931 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9583 GND A3 word161 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9584 a_1766_n134816# A3 a_1370_n134816# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9585 a_974_n131408# A6 a_578_n131408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9586 GND A3 word102 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9587 a_974_n63390# A6 a_578_n63390# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9588 a_314_n116072# a_264_n66# a_50_n116072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9589 word910 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9590 a_2030_n113942# A2 a_1766_n113942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9591 a_1634_n44930# a_1584_n66# a_1370_n44930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9592 GND A5 word531 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9593 word476 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9594 a_578_n93494# a_528_n66# a_446_n93494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9595 a_1238_n83412# A5 a_842_n83412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9596 word684 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9597 GND A4 word45 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9598 a_710_n48622# A7 a_314_n48622# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9599 word966 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9600 word907 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9601 a_974_n130982# A6 a_578_n130982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9602 word63 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9603 a_2162_n106842# a_2112_n66# a_1898_n106842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9604 word688 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9605 a_182_n14400# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9606 word156 A0 a_2294_n22352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9607 word254 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9608 a_446_n25902# A8 a_182_n25902# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9609 a_1898_n44078# a_1848_n66# a_1766_n44078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9610 word195 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9611 a_1634_n99742# a_1584_n66# a_1370_n99742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9612 a_842_n142058# a_792_n66# a_578_n142058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9613 a_1370_n2898# a_1320_n66# a_1238_n2898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9614 word486 A0 a_2162_n69212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9615 word464 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9616 GND A3 word368 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9617 a_1502_n74182# A4 a_1238_n74182# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9618 GND A9 word243 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9619 a_314_n145466# a_264_n66# a_50_n145466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9620 word457 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9621 word94 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9622 a_1766_n102866# A3 a_1370_n102866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9623 a_842_n119196# a_792_n66# a_710_n119196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9624 a_1634_n12980# a_1584_n66# a_1370_n12980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9625 a_1238_n29026# A5 a_842_n29026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9626 word708 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9627 a_2294_n28032# A1 a_1898_n28032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9628 a_842_n71200# a_792_n66# a_578_n71200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9629 a_1634_n68218# a_1584_n66# a_1370_n68218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9630 a_2030_n68502# A2 a_1766_n68502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9631 a_974_n78300# A6 a_710_n78300# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9632 word582 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9633 a_2030_n128852# A2 a_1634_n128852# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9634 a_2162_n12554# a_2112_n66# a_1898_n12554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9635 a_2294_n19654# A1 a_2030_n19654# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9636 a_1634_n90654# a_1584_n66# a_1370_n90654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9637 a_710_n16672# A7 a_446_n16672# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9638 GND A6 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9639 word422 A0 a_2162_n60124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9640 a_1106_n117350# a_1056_n66# a_974_n117350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9641 GND A2 word40 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9642 word358 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9643 a_1634_n140354# a_1584_n66# a_1370_n140354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9644 word299 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9645 word31 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9646 GND A5 word84 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9647 word561 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9648 a_1238_n11560# A5 a_842_n11560# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9649 word292 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9650 a_1634_n67792# a_1584_n66# a_1370_n67792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9651 word202 A0 a_2162_n28884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9652 a_2294_n71910# A1 a_2030_n71910# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9653 word360 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9654 GND A9 word77 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9655 a_1634_n117492# a_1584_n66# a_1370_n117492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9656 a_2294_n10566# A1 a_2030_n10566# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9657 word138 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9658 a_1238_n58420# A5 a_974_n58420# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9659 word622 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9660 GND A9 word348 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9661 GND A6 word811 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9662 word199 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9663 a_1766_n126154# A3 a_1370_n126154# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9664 a_974_n114368# A6 a_710_n114368# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9665 a_2162_n41948# a_2112_n66# a_1898_n41948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9666 word339 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9667 a_1634_n36268# a_1584_n66# a_1370_n36268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9668 a_2030_n36552# A2 a_1766_n36552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9669 a_710_n54444# A7 a_314_n54444# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9670 word357 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9671 word872 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9672 word1007 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9673 GND A5 word411 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9674 word497 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9675 a_2162_n121042# a_2112_n66# a_2030_n121042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9676 a_1238_n57994# A5 a_974_n57994# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9677 a_1238_n66372# A5 a_842_n66372# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9678 a_446_n31724# A8 a_182_n31724# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9679 GND A1 word181 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9680 GND A7 word874 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9681 a_1766_n13832# A3 a_1502_n13832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9682 GND A7 word815 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9683 word468 A0 a_2294_n66656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9684 GND A9 word284 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9685 word877 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9686 a_2294_n125302# A1 a_2030_n125302# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9687 word93 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9688 GND A5 word130 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9689 GND A7 word46 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9690 word465 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9691 GND A7 word871 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9692 GND A9 word182 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9693 GND A9 word123 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9694 a_1238_n122604# A5 a_842_n122604# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9695 word500 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9696 a_1634_n74040# a_1584_n66# a_1502_n74040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9697 a_2030_n74324# A2 a_1634_n74324# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9698 word605 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9699 a_2030_n134674# A2 a_1766_n134674# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9700 GND A4 word736 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9701 a_710_n83838# A7 a_446_n83838# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9702 a_1370_n12412# a_1320_n66# a_1238_n12412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9703 word932 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9704 a_2162_n56858# a_2112_n66# a_1898_n56858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9705 a_2162_n65236# a_2112_n66# a_2030_n65236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9706 a_974_n129278# A6 a_578_n129278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9707 word175 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9708 word661 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9709 word670 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9710 word302 A0 a_2162_n43084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9711 a_1370_n108404# a_1320_n66# a_1106_n108404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9712 word711 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9713 word941 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9714 word710 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9715 GND A9 word61 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9716 GND A2 word512 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9717 GND A3 word514 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9718 GND A9 word389 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9719 word240 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9720 a_2294_n54870# A1 a_2030_n54870# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9721 a_2294_n63248# A1 a_1898_n63248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9722 GND A1 word713 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9723 a_1766_n123598# A3 a_1502_n123598# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9724 word717 a_2376_n66# a_2294_n102014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9725 a_710_n51888# A7 a_314_n51888# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9726 a_2030_n42374# A2 a_1634_n42374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9727 GND A5 word452 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9728 word139 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9729 GND A8 word229 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9730 word854 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9731 GND A1 word984 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9732 a_1238_n137514# A5 a_842_n137514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9733 word707 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9734 word912 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9735 a_446_n15110# A8 a_182_n15110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9736 GND A7 word82 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9737 a_2030_n89234# A2 a_1766_n89234# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9738 a_710_n113232# A7 a_314_n113232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9739 GND A4 word841 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9740 GND A1 word281 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9741 a_1370_n27322# a_1320_n66# a_1106_n27322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9742 word686 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9743 GND A8 word127 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9744 GND A0 word822 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9745 a_446_n84406# A8 a_50_n84406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9746 a_1766_n66514# A3 a_1370_n66514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9747 word716 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9748 word626 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9749 a_446_n23062# A8 a_182_n23062# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9750 GND A6 word56 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9751 a_446_n14684# A8 a_182_n14684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9752 word75 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9753 word438 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9754 a_1106_n5028# a_1056_n66# a_974_n5028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9755 GND A2 word129 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9756 word848 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9757 GND A9 word164 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9758 GND A1 word920 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9759 a_2030_n80146# A2 a_1766_n80146# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9760 word757 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9761 GND A4 word777 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9762 a_578_n142342# a_528_n66# a_314_n142342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9763 a_578_n133964# a_528_n66# a_314_n133964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9764 a_2030_n71768# A2 a_1634_n71768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9765 GND A5 word659 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9766 a_2294_n108262# A1 a_2030_n108262# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9767 a_2294_n78158# A1 a_1898_n78158# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9768 GND A2 word617 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9769 GND A6 word957 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9770 a_2162_n71058# a_2112_n66# a_2030_n71058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9771 word345 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9772 a_446_n102156# A8 a_50_n102156# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9773 a_974_n135100# A6 a_578_n135100# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9774 a_710_n75176# A7 a_446_n75176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9775 a_2030_n57284# A2 a_1766_n57284# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9776 word485 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9777 word763 a_2376_n66# a_2162_n108546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9778 word921 a_2376_n66# a_2294_n130982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9779 word461 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9780 a_2162_n133396# a_2112_n66# a_2030_n133396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9781 word824 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9782 word727 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9783 word391 a_2376_n66# a_2162_n55722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9784 a_578_n102440# a_528_n66# a_446_n102440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9785 a_1766_n95908# A3 a_1502_n95908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9786 word765 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9787 a_50_n104712# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9788 a_2162_n48196# a_2112_n66# a_2030_n48196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9789 a_710_n119764# A7 a_314_n119764# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9790 a_1766_n34564# A3 a_1370_n34564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9791 word614 A0 a_2162_n87388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9792 GND A9 word430 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9793 GND A5 word729 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9794 word1023 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9795 a_1502_n114510# A4 a_1106_n114510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9796 a_1106_n15536# a_1056_n66# a_842_n15536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9797 a_446_n99316# A8 a_50_n99316# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9798 word550 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9799 a_2294_n137656# A1 a_2030_n137656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9800 a_446_n29594# A8 a_182_n29594# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9801 word239 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9802 a_1502_n342# A4 a_1238_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9803 GND A1 word52 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9804 word953 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9805 GND A2 word451 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9806 GND A9 word269 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9807 GND A1 word105 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9808 GND A2 word392 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9809 a_2030_n86678# A2 a_1766_n86678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9810 a_710_n9714# A7 a_446_n9714# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9811 GND A8 word7 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9812 a_710_n110676# A7 a_314_n110676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9813 a_1370_n143620# a_1320_n66# a_1106_n143620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9814 GND A0 word922 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9815 a_842_n16814# a_792_n66# a_710_n16814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9816 GND A8 word168 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9817 word1019 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9818 a_446_n90228# A8 a_50_n90228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9819 GND A8 word109 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9820 GND A1 word593 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9821 a_446_n81850# A8 a_50_n81850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9822 a_1766_n63958# A3 a_1502_n63958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9823 a_446_n108688# A8 a_50_n108688# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9824 GND A1 word161 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9825 GND A6 word38 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9826 a_1106_n53308# a_1056_n66# a_842_n53308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9827 GND A7 word795 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9828 GND A8 word656 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9829 GND A2 word170 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9830 a_1106_n44930# a_1056_n66# a_974_n44930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9831 GND A6 word293 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9832 GND A8 word597 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9833 a_50_n119622# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9834 GND A8 word726 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9835 word57 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9836 a_1502_n129420# A4 a_1238_n129420# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9837 GND A5 word834 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9838 a_974_n23204# A6 a_578_n23204# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9839 GND A2 word658 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9840 GND A6 word132 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9841 GND A6 word191 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9842 a_1238_n111386# A5 a_974_n111386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9843 GND A3 word804 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9844 GND A1 word800 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9845 GND A2 word226 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9846 a_1106_n52882# a_1056_n66# a_842_n52882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9847 a_50_n75602# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9848 word344 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9849 a_1370_n62538# a_1320_n66# a_1106_n62538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9850 word745 a_2376_n66# a_2294_n105990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9851 word1000 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9852 a_1106_n99742# a_1056_n66# a_974_n99742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9853 a_1370_n111670# a_1320_n66# a_1238_n111670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9854 a_50_n110534# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9855 a_1502_n137372# A4 a_1238_n137372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9856 a_1502_n128994# A4 a_1238_n128994# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9857 a_710_n125586# A7 a_314_n125586# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9858 GND A1 word368 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9859 a_1370_n39676# a_1320_n66# a_1238_n39676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9860 a_1370_n48054# a_1320_n66# a_1238_n48054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9861 GND A0 word968 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9862 GND A7 word558 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9863 a_446_n96760# A8 a_50_n96760# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9864 a_1766_n87246# A3 a_1502_n87246# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9865 word122 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9866 GND A7 word126 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9867 word271 a_2376_n66# a_2162_n38682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9868 a_2294_n143478# A1 a_2030_n143478# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9869 GND A2 word275 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9870 a_1106_n59840# a_1056_n66# a_974_n59840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9871 word994 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9872 GND A6 word398 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9873 a_1106_n90654# a_1056_n66# a_842_n90654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9874 word935 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9875 GND A8 word702 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9876 a_1238_n140780# A5 a_842_n140780# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9877 GND A2 word433 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9878 a_2030_n92500# A2 a_1634_n92500# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9879 GND A4 word864 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9880 a_974_n38114# A6 a_710_n38114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9881 GND A5 word21 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9882 word117 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9883 a_842_n31014# a_792_n66# a_578_n31014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9884 a_1370_n30588# a_1320_n66# a_1238_n30588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9885 word639 a_2376_n66# a_2162_n90938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9886 GND A1 word964 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9887 GND A2 word962 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9888 GND A8 word150 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9889 word833 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9890 word909 a_2376_n66# a_2294_n129278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9891 a_314_n41522# a_264_n66# a_182_n41522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9892 word607 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9893 GND A0 word802 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9894 a_1898_n24908# a_1848_n66# a_1634_n24908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9895 word537 a_2376_n66# a_2294_n76454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9896 GND A8 word638 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9897 a_1370_n126580# a_1320_n66# a_1106_n126580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9898 a_446_n2046# A8 a_182_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9899 a_50_n125444# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9900 a_1898_n7726# a_1848_n66# a_1766_n7726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9901 GND A0 word456 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9902 GND A1 word473 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9903 GND A7 word333 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9904 a_446_n73188# A8 a_50_n73188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9905 a_1766_n55296# A3 a_1502_n55296# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9906 word381 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9907 word322 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9908 a_974_n20648# A6 a_578_n20648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9909 a_1106_n36268# a_1056_n66# a_842_n36268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9910 a_578_n28316# a_528_n66# a_446_n28316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9911 GND A6 word173 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9912 a_842_n108404# a_792_n66# a_578_n108404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9913 a_578_n19938# a_528_n66# a_446_n19938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9914 word845 a_2376_n66# a_2294_n120190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9915 a_50_n81424# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9916 GND A3 word131 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9917 GND A0 word234 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9918 a_578_n97612# a_528_n66# a_446_n97612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9919 GND A2 word538 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9920 a_1502_n143194# A4 a_1106_n143194# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9921 GND A2 word737 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9922 GND A4 word969 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9923 a_314_n70916# a_264_n66# a_182_n70916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9924 GND A4 word227 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9925 a_1370_n45498# a_1320_n66# a_1106_n45498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9926 GND A7 word540 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9927 GND A7 word599 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9928 word798 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9929 GND A1 word680 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9930 a_1766_n84690# A3 a_1370_n84690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9931 a_182_n18518# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9932 a_314_n56432# a_264_n66# a_182_n56432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9933 word978 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9934 a_182_n40954# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9935 a_314_n111102# a_264_n66# a_50_n111102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9936 a_578_n57710# a_528_n66# a_314_n57710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9937 a_1898_n39818# a_1848_n66# a_1766_n39818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9938 GND A6 word439 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9939 word441 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9940 a_446_n8578# A8 a_182_n8578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9941 word48 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9942 a_446_n88098# A8 a_50_n88098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9943 word942 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9944 GND A4 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9945 a_1502_n69922# A4 a_1106_n69922# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9946 GND A5 word980 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9947 word486 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9948 word946 A0 a_2162_n134532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9949 word158 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9950 word931 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9951 GND A2 word1003 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9952 GND A3 word950 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9953 GND A6 word278 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9954 word739 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9955 a_578_n65662# a_528_n66# a_314_n65662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9956 GND A4 word493 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9957 word653 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9958 a_50_n96334# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9959 a_50_n87956# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9960 a_842_n66940# a_792_n66# a_578_n66940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9961 word160 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9962 word1005 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9963 a_1634_n9146# a_1584_n66# a_1370_n9146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9964 a_1898_n30730# a_1848_n66# a_1766_n30730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9965 word519 a_2376_n66# a_2162_n73898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9966 word646 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9967 word724 A0 a_2294_n103008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9968 a_50_n131266# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9969 GND A0 word280 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9970 word370 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9971 word551 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9972 GND A2 word842 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9973 a_50_n122888# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9974 GND A4 word332 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9975 a_1502_n60834# A4 a_1106_n60834# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9976 a_1106_n143904# a_1056_n66# a_842_n143904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9977 word422 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9978 word363 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9979 a_1106_n42090# a_1056_n66# a_974_n42090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9980 word903 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9981 a_578_n34138# a_528_n66# a_446_n34138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9982 GND A6 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9983 word216 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9984 a_842_n105848# a_792_n66# a_578_n105848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9985 a_578_n25760# a_528_n66# a_446_n25760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9986 word15 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9987 GND A3 word231 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9988 word209 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9989 a_182_n64242# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9990 a_974_n73330# A6 a_710_n73330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9991 a_314_n126012# a_264_n66# a_50_n126012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9992 a_182_n55864# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9993 a_1502_n37972# A4 a_1238_n37972# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9994 a_314_n117634# a_264_n66# a_50_n117634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X9995 GND A6 word544 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X9996 word261 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9997 a_2294_n1478# A1 a_2030_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9998 a_710_n11702# A7 a_446_n11702# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X9999 a_1502_n6022# A4 a_1106_n6022# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10000 word706 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10001 GND A2 word778 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10002 word263 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10003 a_842_n34990# a_792_n66# a_578_n34990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10004 a_1634_n62822# a_1584_n66# a_1370_n62822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10005 a_974_n81282# A6 a_710_n81282# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10006 word977 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10007 word780 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10008 a_182_n6164# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10009 GND A0 word114 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10010 a_1370_n98180# a_1320_n66# a_1106_n98180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10011 word1002 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10012 a_182_n24340# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10013 a_314_n62254# a_264_n66# a_182_n62254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10014 word145 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10015 a_314_n53876# a_264_n66# a_182_n53876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10016 GND A4 word107 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10017 word162 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10018 word103 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10019 word534 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10020 word683 a_2376_n66# a_2162_n97186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10021 a_842_n143620# a_792_n66# a_578_n143620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10022 a_50_n137798# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10023 GND A3 word20 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10024 word475 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10025 a_1502_n84122# A4 a_1238_n84122# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10026 GND A0 word602 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10027 word770 A0 a_2162_n109540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10028 word62 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10029 word96 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10030 word928 A0 a_2294_n131976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10031 word755 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10032 word468 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10033 a_182_n32292# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10034 a_314_n39392# a_264_n66# a_182_n39392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10035 a_974_n41380# A6 a_710_n41380# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10036 GND A6 word319 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10037 word10 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10038 a_578_n71484# a_528_n66# a_314_n71484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10039 a_50_n93778# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10040 GND A3 word277 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10041 word826 A0 a_2162_n117492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10042 word470 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10043 a_1634_n6590# a_1584_n66# a_1502_n6590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10044 GND A0 word380 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10045 a_3028_164# A0 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X10046 word592 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10047 word811 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10048 word752 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10049 GND A2 word883 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10050 a_1634_n30872# a_1584_n66# a_1370_n30872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10051 word301 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10052 word533 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10053 a_50_n79294# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10054 a_842_n49900# a_792_n66# a_710_n49900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10055 word491 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10056 a_974_n96192# A6 a_578_n96192# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10057 word362 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10058 word526 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10059 word631 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10060 word885 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10061 a_842_n120048# a_792_n66# a_710_n120048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10062 a_182_n39250# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10063 a_1898_n13690# a_1848_n66# a_1634_n13690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10064 word250 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10065 word309 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10066 a_314_n68786# a_264_n66# a_182_n68786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10067 a_182_n70064# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10068 GND A3 word213 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10069 word272 A0 a_2294_n38824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10070 a_1502_n52172# A4 a_1106_n52172# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10071 a_1106_n135242# a_1056_n66# a_974_n135242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10072 a_182_n61686# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10073 word267 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10074 a_314_n123456# a_264_n66# a_50_n123456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10075 word302 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10076 a_1106_n126864# a_1056_n66# a_842_n126864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10077 word79 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10078 GND A3 word484 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10079 a_1898_n82986# a_1848_n66# a_1766_n82986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10080 GND A5 word151 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10081 GND A6 word822 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10082 a_1766_n127716# A3 a_1502_n127716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10083 a_974_n115930# A6 a_710_n115930# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10084 word245 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10085 a_1634_n37830# a_1584_n66# a_1502_n37830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10086 a_974_n56290# A6 a_578_n56290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10087 word567 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10088 word1018 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10089 a_1238_n67934# A5 a_842_n67934# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10090 a_1238_n76312# A5 a_974_n76312# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10091 GND A4 word580 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10092 a_2162_n122604# a_2112_n66# a_1898_n122604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10093 word736 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10094 a_2162_n37404# a_2112_n66# a_1898_n37404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10095 word719 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10096 word697 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10097 word44 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10098 word474 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10099 GND A0 word34 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10100 word106 A0 a_2162_n15252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10101 GND A4 word419 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10102 word509 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10103 word204 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10104 a_1898_n135952# a_1848_n66# a_1634_n135952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10105 a_1370_n4176# a_1320_n66# a_1238_n4176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10106 a_446_n18802# A8 a_182_n18802# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10107 a_842_n126580# a_792_n66# a_710_n126580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10108 GND A9 word193 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10109 GND A3 word259 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10110 a_314_n138366# a_264_n66# a_50_n138366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10111 a_2030_n144614# A2 a_1634_n144614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10112 a_2294_n35416# A1 a_2030_n35416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10113 a_314_n129988# a_264_n66# a_50_n129988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10114 word692 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10115 GND A6 word690 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10116 a_1502_n9998# A4 a_1238_n9998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10117 word125 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10118 GND A5 word256 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10119 word633 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10120 word852 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10121 word717 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10122 a_1898_n104428# a_1848_n66# a_1634_n104428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10123 word591 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10124 word350 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10125 a_842_n64100# a_792_n66# a_578_n64100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10126 word140 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10127 a_1634_n83554# a_1584_n66# a_1502_n83554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10128 a_2162_n137514# a_2112_n66# a_1898_n137514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10129 GND A2 word49 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10130 word372 A0 a_2294_n53024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10131 GND A4 word685 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10132 GND A3 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10133 a_1106_n141064# a_1056_n66# a_842_n141064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10134 a_1634_n133254# a_1584_n66# a_1502_n133254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10135 word781 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10136 a_314_n120900# a_264_n66# a_50_n120900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10137 a_1106_n132686# a_1056_n66# a_974_n132686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10138 a_1634_n124876# a_1584_n66# a_1502_n124876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10139 word674 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10140 word242 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10141 GND A6 word922 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10142 a_1502_n96476# A4 a_1106_n96476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10143 a_2030_n121042# A2 a_1766_n121042# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10144 a_974_n130130# A6 a_578_n130130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10145 a_1634_n52030# a_1584_n66# a_1502_n52030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10146 a_2030_n112664# A2 a_1634_n112664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10147 GND A5 word463 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10148 GND A5 word522 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10149 a_1238_n73756# A5 a_974_n73756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10150 a_1238_n82134# A5 a_842_n82134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10151 a_1766_n119054# A3 a_1502_n119054# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10152 a_2162_n43226# a_2112_n66# a_1898_n43226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10153 GND A9 word456 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10154 a_1634_n29168# a_1584_n66# a_1502_n29168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10155 a_710_n47344# A7 a_314_n47344# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10156 GND A8 word36 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10157 word366 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10158 word957 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10159 a_710_n38966# A7 a_314_n38966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10160 word447 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10161 word515 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10162 a_2162_n105564# a_2112_n66# a_1898_n105564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10163 word763 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10164 a_1898_n119338# a_1848_n66# a_1766_n119338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10165 word88 A0 a_2294_n12696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10166 a_446_n33002# A8 a_182_n33002# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10167 a_1898_n141774# a_1848_n66# a_1766_n141774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10168 a_446_n24624# A8 a_182_n24624# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10169 GND A1 word17 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10170 word508 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10171 GND A7 word824 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10172 word418 A0 a_2162_n59556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10173 GND A9 word234 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10174 GND A3 word359 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10175 a_314_n144188# a_264_n66# a_50_n144188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10176 word827 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10177 word85 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10178 a_2294_n41238# A1 a_2030_n41238# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10179 word576 A0 a_2294_n81992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10180 a_578_n143904# a_528_n66# a_314_n143904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10181 a_1634_n20080# a_1584_n66# a_1502_n20080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10182 word225 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10183 word571 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10184 GND A3 word689 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10185 a_2294_n109824# A1 a_1898_n109824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10186 a_2030_n11986# A2 a_1766_n11986# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10187 GND A3 word630 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10188 a_842_n9572# a_792_n66# a_710_n9572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10189 a_1238_n19370# A5 a_974_n19370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10190 a_2162_n72620# a_2112_n66# a_1898_n72620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10191 GND A8 word74 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10192 a_2294_n79720# A1 a_2030_n79720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10193 GND A1 word829 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10194 a_710_n85116# A7 a_446_n85116# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10195 a_446_n103718# A8 a_50_n103718# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10196 word555 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10197 GND A7 word821 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10198 a_1898_n110250# a_1848_n66# a_1766_n110250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10199 a_2162_n11276# a_2112_n66# a_1898_n11276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10200 a_2294_n18376# A1 a_2030_n18376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10201 a_710_n76738# A7 a_446_n76738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10202 a_2030_n67224# A2 a_1634_n67224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10203 a_2030_n127574# A2 a_1766_n127574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10204 a_1634_n80998# a_1584_n66# a_1370_n80998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10205 word970 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10206 word991 a_2376_n66# a_2162_n140922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10207 a_710_n15394# A7 a_446_n15394# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10208 word354 A0 a_2162_n50468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10209 word290 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10210 a_2294_n87672# A1 a_2030_n87672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10211 word471 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10212 a_2162_n80572# a_2112_n66# a_1898_n80572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10213 a_2294_n100736# A1 a_1898_n100736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10214 word684 A0 a_2294_n97328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10215 word891 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10216 word613 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10217 word554 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10218 GND A3 word464 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10219 GND A9 word339 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10220 GND A6 word802 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10221 GND A9 word280 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10222 a_1502_n132402# A4 a_1106_n132402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10223 a_974_n113090# A6 a_710_n113090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10224 GND A9 word497 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10225 a_1766_n116498# A3 a_1370_n116498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10226 a_710_n120616# A7 a_314_n120616# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10227 a_710_n53166# A7 a_314_n53166# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10228 GND A8 word18 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10229 a_710_n44788# A7 a_314_n44788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10230 a_1370_n34706# a_1320_n66# a_1106_n34706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10231 GND A5 word402 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10232 a_1238_n65094# A5 a_842_n65094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10233 GND A8 word179 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10234 a_2162_n87530# a_2112_n66# a_1898_n87530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10235 word745 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10236 a_2162_n111386# a_2112_n66# a_1898_n111386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10237 GND A7 word91 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10238 a_2162_n26186# a_2112_n66# a_1898_n26186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10239 a_446_n30446# A8 a_182_n30446# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10240 a_1766_n12554# A3 a_1370_n12554# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10241 GND A1 word172 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10242 GND A7 word865 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10243 GND A9 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10244 GND A8 word667 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10245 GND A0 word772 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10246 word400 A0 a_2294_n57000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10247 a_446_n77306# A8 a_50_n77306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10248 word395 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10249 a_1766_n59414# A3 a_1502_n59414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10250 a_2162_n95482# a_2112_n66# a_1898_n95482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10251 GND A8 word737 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10252 a_2294_n124024# A1 a_2030_n124024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10253 a_2294_n115646# A1 a_1898_n115646# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10254 GND A7 word37 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10255 word798 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10256 GND A1 word929 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10257 a_1238_n121326# A5 a_842_n121326# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10258 GND A2 word296 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10259 a_1106_n62822# a_1056_n66# a_974_n62822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10260 GND A9 word114 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10261 a_578_n135242# a_528_n66# a_314_n135242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10262 a_1238_n112948# A5 a_974_n112948# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10263 a_2294_n24198# A1 a_2030_n24198# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10264 a_2030_n73046# A2 a_1766_n73046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10265 a_710_n82560# A7 a_446_n82560# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10266 a_1502_n100452# A4 a_1238_n100452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10267 GND A5 word668 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10268 a_2030_n133396# A2 a_1634_n133396# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10269 word815 a_2376_n66# a_2162_n115930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10270 word572 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10271 a_1238_n94488# A5 a_974_n94488# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10272 word923 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10273 a_2162_n140780# a_2112_n66# a_1898_n140780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10274 a_1370_n121610# a_1320_n66# a_1238_n121610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10275 GND A7 word298 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10276 GND A0 word708 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10277 GND A1 word768 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10278 a_974_n4318# A6 a_710_n4318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10279 a_1766_n50326# A3 a_1502_n50326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10280 a_2162_n55580# a_2112_n66# a_1898_n55580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10281 a_2294_n93494# A1 a_2030_n93494# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10282 GND A9 word55 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10283 a_2162_n1762# a_2112_n66# a_2030_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10284 a_1766_n41948# A3 a_1502_n41948# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10285 GND A3 word871 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10286 a_1370_n49616# a_1320_n66# a_1238_n49616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10287 word871 a_2376_n66# a_2162_n123882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10288 a_1106_n22920# a_1056_n66# a_974_n22920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10289 word411 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10290 a_1370_n107126# a_1320_n66# a_1106_n107126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10291 word341 a_2376_n66# a_2294_n48622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10292 a_1766_n88808# A3 a_1370_n88808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10293 GND A1 word277 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10294 a_1766_n27464# A3 a_1502_n27464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10295 a_974_n3892# A6 a_710_n3892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10296 GND A2 word562 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10297 word1005 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10298 GND A9 word380 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10299 GND A9 word52 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10300 GND A1 word704 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10301 GND A4 word993 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10302 word973 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10303 GND A4 word934 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10304 a_2030_n41096# A2 a_1766_n41096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10305 a_578_n103292# a_528_n66# a_446_n103292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10306 word189 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10307 a_1370_n40528# a_1320_n66# a_1238_n40528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10308 word845 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10309 GND A8 word220 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10310 word903 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10311 GND A3 word979 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10312 GND A2 word401 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10313 a_1106_n77732# a_1056_n66# a_974_n77732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10314 word979 a_2376_n66# a_2162_n139218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10315 a_1238_n127858# A5 a_974_n127858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10316 GND A4 word832 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10317 a_1502_n115362# A4 a_1106_n115362# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10318 GND A7 word73 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10319 GND A4 word773 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10320 GND A1 word213 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10321 word884 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10322 a_1370_n17666# a_1320_n66# a_1106_n17666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10323 a_1370_n26044# a_1320_n66# a_1106_n26044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10324 word500 A0 a_2294_n71200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10325 word618 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10326 word969 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10327 GND A0 word872 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10328 a_446_n3608# A8 a_182_n3608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10329 a_446_n74750# A8 a_50_n74750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10330 a_446_n83128# A8 a_50_n83128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10331 GND A1 word484 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10332 GND A3 word976 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10333 GND A2 word120 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10334 GND A8 word606 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10335 GND A3 word915 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10336 GND A7 word19 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10337 word780 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10338 GND A8 word547 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10339 a_1370_n144472# a_1320_n66# a_1106_n144472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10340 word915 a_2376_n66# a_2162_n130130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10341 a_578_n141064# a_528_n66# a_314_n141064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10342 GND A4 word709 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10343 a_578_n132686# a_528_n66# a_314_n132686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10344 GND A5 word650 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10345 word700 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10346 GND A9 word485 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10347 GND A2 word608 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10348 GND A1 word809 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10349 GND A3 word754 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10350 GND A2 word176 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10351 a_1238_n104286# A5 a_842_n104286# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10352 GND A7 word610 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10353 a_1370_n104570# a_1320_n66# a_1238_n104570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10354 a_50_n103434# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10355 a_710_n118486# A7 a_314_n118486# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10356 GND A4 word136 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10357 GND A5 word720 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10358 a_1106_n14258# a_1056_n66# a_842_n14258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10359 a_446_n98038# A8 a_50_n98038# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10360 a_446_n89660# A8 a_50_n89660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10361 a_2294_n128000# A1 a_1898_n128000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10362 word944 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10363 word885 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10364 GND A4 word873 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10365 GND A5 word776 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10366 a_710_n8436# A7 a_446_n8436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10367 a_2030_n85400# A2 a_1634_n85400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10368 GND A4 word814 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10369 word925 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10370 GND A4 word72 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10371 GND A0 word854 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10372 a_842_n15536# a_792_n66# a_710_n15536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10373 a_50_n141206# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10374 GND A8 word100 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10375 word589 a_2376_n66# a_2294_n83838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10376 GND A2 word912 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10377 a_1238_n119196# A5 a_842_n119196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10378 a_50_n132828# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10379 a_1766_n71058# A3 a_1370_n71058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10380 GND A1 word525 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10381 GND A1 word584 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10382 word157 a_2376_n66# a_2294_n22494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10383 word806 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10384 GND A0 word76 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10385 a_1106_n52030# a_1056_n66# a_842_n52030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10386 word557 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10387 word823 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10388 GND A6 word284 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10389 word487 a_2376_n66# a_2162_n69354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10390 a_842_n84832# a_792_n66# a_710_n84832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10391 GND A8 word647 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10392 GND A8 word588 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10393 word764 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10394 a_50_n118344# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10395 a_1898_n9004# a_1848_n66# a_1634_n9004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10396 a_1898_n17808# a_1848_n66# a_1634_n17808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10397 word1019 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10398 word846 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10399 a_50_n109966# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10400 word279 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10401 a_1766_n48196# A3 a_1370_n48196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10402 GND A0 word406 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10403 word496 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10404 word787 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10405 a_182_n65804# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10406 word331 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10407 word19 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10408 word272 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10409 a_1634_n1620# a_1584_n66# a_1502_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10410 GND A6 word182 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10411 GND A2 word649 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10412 GND A2 word848 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10413 word795 a_2376_n66# a_2162_n113090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10414 a_50_n74324# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10415 a_842_n53308# a_792_n66# a_710_n53308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10416 a_974_n91222# A6 a_578_n91222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10417 a_1106_n98464# a_1056_n66# a_974_n98464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10418 GND A0 word184 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10419 word423 a_2376_n66# a_2162_n60266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10420 GND A2 word488 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10421 GND A2 word746 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10422 a_182_n7726# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10423 a_50_n100878# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10424 word215 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10425 a_314_n63816# a_264_n66# a_182_n63816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10426 word2 A0 a_2162_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10427 GND A1 word300 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10428 GND A7 word549 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10429 GND A0 word900 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10430 GND A0 word672 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10431 GND A1 word689 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10432 word748 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10433 a_842_n52882# a_792_n66# a_710_n52882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10434 a_974_n59982# A6 a_578_n59982# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10435 a_1766_n77590# A3 a_1502_n77590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10436 a_2294_n142200# A1 a_2030_n142200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10437 word998 A0 a_2162_n141916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10438 word113 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10439 a_182_n42232# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10440 a_314_n49332# a_264_n66# a_182_n49332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10441 a_182_n33854# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10442 a_1502_n15962# A4 a_1106_n15962# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10443 GND A6 word389 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10444 word391 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10445 word985 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10446 a_1898_n63532# a_1848_n66# a_1634_n63532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10447 a_1106_n80998# a_1056_n66# a_974_n80998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10448 word951 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10449 word601 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10450 word896 A0 a_2294_n127432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10451 a_710_n5880# A7 a_446_n5880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10452 a_974_n484# A6 a_710_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10453 a_842_n12980# a_792_n66# a_710_n12980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10454 word13 a_2376_n66# a_2294_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10455 word108 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10456 word881 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10457 word822 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10458 GND A2 word953 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10459 a_1634_n40812# a_1584_n66# a_1370_n40812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10460 word603 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10461 word662 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10462 a_50_n89234# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10463 a_578_n58562# a_528_n66# a_314_n58562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10464 GND A4 word384 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10465 a_1370_n76170# a_1320_n66# a_1238_n76170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10466 a_314_n40244# a_264_n66# a_182_n40244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10467 a_842_n68218# a_792_n66# a_578_n68218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10468 a_842_n90654# a_792_n66# a_710_n90654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10469 word596 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10470 a_974_n97754# A6 a_578_n97754# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10471 a_50_n124166# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10472 a_1898_n6448# a_1848_n66# a_1634_n6448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10473 a_1898_n23630# a_1848_n66# a_1766_n23630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10474 word379 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10475 word469 a_2376_n66# a_2294_n66798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10476 GND A0 word506 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10477 a_842_n121610# a_792_n66# a_710_n121610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10478 a_50_n115788# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10479 GND A1 word464 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10480 a_182_n71626# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10481 GND A6 word655 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10482 word372 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10483 word313 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10484 a_182_n10282# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10485 a_842_n107126# a_792_n66# a_578_n107126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10486 a_1898_n92926# a_1848_n66# a_1634_n92926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10487 a_578_n18660# a_528_n66# a_446_n18660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10488 a_578_n27038# a_528_n66# a_446_n27038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10489 GND A6 word164 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10490 a_842_n67792# a_792_n66# a_578_n67792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10491 word166 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10492 word726 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10493 a_1898_n31582# a_1848_n66# a_1634_n31582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10494 a_182_n48764# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10495 a_182_n57142# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10496 a_50_n80146# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10497 word374 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10498 word376 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10499 a_578_n96334# a_528_n66# a_446_n96334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10500 a_1898_n78442# a_1848_n66# a_1766_n78442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10501 GND A2 word728 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10502 GND A6 word652 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10503 GND A4 word65 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10504 GND A0 word1000 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10505 a_1766_n7158# A3 a_1370_n7158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10506 word59 a_2376_n66# a_2162_n8578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10507 a_842_n27890# a_792_n66# a_578_n27890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10508 a_842_n36268# a_792_n66# a_578_n36268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10509 a_974_n74182# A6 a_710_n74182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10510 word336 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10511 a_974_n133822# A6 a_578_n133822# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10512 word789 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10513 GND A4 word548 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10514 a_1502_n91506# A4 a_1238_n91506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10515 a_182_n17240# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10516 word95 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10517 word154 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10518 GND A4 word489 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10519 word952 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10520 a_314_n46776# a_264_n66# a_182_n46776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10521 a_314_n55154# a_264_n66# a_182_n55154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10522 GND A2 word11 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10523 GND A6 word430 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10524 a_1106_n104854# a_1056_n66# a_842_n104854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10525 word701 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10526 word432 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10527 a_842_n136520# a_792_n66# a_578_n136520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10528 a_50_n139076# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10529 a_1898_n38540# a_1848_n66# a_1634_n38540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10530 a_446_n7300# A8 a_182_n7300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10531 a_1898_n60976# a_1848_n66# a_1634_n60976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10532 GND A0 word552 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10533 a_1502_n68644# A4 a_1106_n68644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10534 a_314_n139928# a_264_n66# a_50_n139928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10535 a_1766_n105706# A3 a_1502_n105706# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10536 word878 A0 a_2162_n124876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10537 a_182_n25192# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10538 word418 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10539 a_1634_n15820# a_1584_n66# a_1502_n15820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10540 word149 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10541 GND A6 word269 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10542 word922 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10543 word863 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10544 GND A2 word994 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10545 word644 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10546 a_842_n144472# a_792_n66# a_578_n144472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10547 a_50_n95056# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10548 a_578_n64384# a_528_n66# a_314_n64384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10549 a_1238_n45924# A5 a_842_n45924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10550 a_1898_n46492# a_1848_n66# a_1766_n46492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10551 GND A4 word425 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10552 a_50_n86678# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10553 word420 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10554 word479 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10555 word210 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10556 a_2294_n9288# A1 a_2030_n9288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10557 GND A0 word330 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10558 word637 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10559 word111 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10560 word761 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10561 GND A2 word833 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10562 a_1502_n37120# A4 a_1238_n37120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10563 word251 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10564 word542 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10565 GND A4 word264 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10566 GND A4 word323 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10567 a_1106_n142626# a_1056_n66# a_842_n142626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10568 a_314_n130840# a_264_n66# a_50_n130840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10569 word354 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10570 word476 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10571 word894 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10572 word312 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10573 a_842_n104570# a_792_n66# a_578_n104570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10574 GND A3 word163 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10575 GND A7 word786 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10576 a_182_n54586# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10577 a_1502_n36694# A4 a_1238_n36694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10578 a_314_n116356# a_264_n66# a_50_n116356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10579 a_2294_n13406# A1 a_1898_n13406# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10580 GND A6 word535 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10581 a_710_n10424# A7 a_446_n10424# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10582 a_578_n93778# a_528_n66# a_446_n93778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10583 a_1898_n75886# a_1848_n66# a_1766_n75886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10584 word688 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10585 GND A6 word831 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10586 GND A6 word772 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10587 a_1238_n22352# A5 a_974_n22352# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10588 a_974_n117208# A6 a_710_n117208# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10589 word254 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10590 a_2294_n82702# A1 a_1898_n82702# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10591 a_710_n48906# A7 a_314_n48906# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10592 word377 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10593 word517 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10594 word968 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10595 word991 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10596 a_314_n52598# a_264_n66# a_182_n52598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10597 word158 A0 a_2162_n22636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10598 a_1634_n111244# a_1584_n66# a_1502_n111244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10599 word94 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10600 a_974_n116782# A6 a_710_n116782# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10601 a_1634_n38682# a_1584_n66# a_1502_n38682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10602 GND A3 word370 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10603 a_1502_n74466# A4 a_1238_n74466# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10604 word646 A0 a_2162_n91932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10605 a_1766_n111528# A3 a_1370_n111528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10606 word582 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10607 word459 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10608 word400 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10609 a_2030_n21926# A2 a_1634_n21926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10610 word417 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10611 a_1238_n29310# A5 a_842_n29310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10612 a_842_n119480# a_792_n66# a_710_n119480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10613 GND A7 word891 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10614 a_182_n69496# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10615 a_50_n92500# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10616 GND A3 word209 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10617 GND A9 word301 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10618 a_2294_n50752# A1 a_1898_n50752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10619 word211 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10620 a_1634_n90938# a_1584_n66# a_1370_n90938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10621 word802 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10622 a_710_n16956# A7 a_446_n16956# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10623 GND A5 word206 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10624 word351 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10625 word424 A0 a_2294_n60408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10626 a_1238_n37262# A5 a_974_n37262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10627 a_1634_n140638# a_1584_n66# a_1370_n140638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10628 a_1238_n28884# A5 a_842_n28884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10629 word482 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10630 a_1634_n76454# a_1584_n66# a_1370_n76454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10631 word294 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10632 word353 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10633 word731 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10634 GND A9 word79 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10635 GND A3 word145 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10636 a_314_n122178# a_264_n66# a_50_n122178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10637 a_1106_n125586# a_1056_n66# a_842_n125586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10638 word199 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10639 a_314_n113800# a_264_n66# a_50_n113800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10640 word624 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10641 a_1634_n117776# a_1584_n66# a_1370_n117776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10642 GND A3 word534 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10643 a_1502_n2188# A4 a_1238_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10644 GND A5 word142 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10645 GND A6 word813 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10646 GND A5 word83 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10647 a_2162_n50610# a_2112_n66# a_2030_n50610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10648 a_2294_n57710# A1 a_1898_n57710# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10649 word295 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10650 word687 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10651 a_2030_n36836# A2 a_1766_n36836# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10652 GND A5 word472 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10653 word1009 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10654 GND A9 word76 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10655 GND A5 word413 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10656 a_1238_n75034# A5 a_974_n75034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10657 word874 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10658 a_1238_n66656# A5 a_842_n66656# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10659 word727 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10660 a_2162_n112948# a_2112_n66# a_2030_n112948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10661 GND A9 word406 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10662 a_2162_n27748# a_2112_n66# a_2030_n27748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10663 a_2294_n65662# A1 a_1898_n65662# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10664 GND A9 word17 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10665 word397 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10666 word470 A0 a_2162_n66940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10667 word500 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10668 word871 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10669 a_1898_n143052# a_1848_n66# a_1634_n143052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10670 a_446_n17524# A8 a_182_n17524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10671 GND A3 word309 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10672 GND A9 word184 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10673 a_314_n137088# a_264_n66# a_50_n137088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10674 word526 A0 a_2162_n74892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10675 GND A9 word125 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10676 a_2030_n143336# A2 a_1766_n143336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10677 a_578_n136804# a_528_n66# a_314_n136804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10678 word32 A0 a_2294_n4744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10679 a_2294_n25760# A1 a_1898_n25760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10680 word683 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10681 word175 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10682 word993 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10683 word934 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10684 a_1898_n103150# a_1848_n66# a_1766_n103150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10685 GND A7 word771 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10686 a_1106_n7442# a_1056_n66# a_974_n7442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10687 word81 a_2376_n66# a_2294_n11702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10688 a_710_n78016# A7 a_446_n78016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10689 GND A1 word996 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10690 word663 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10691 word979 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10692 word941 a_2376_n66# a_2294_n133822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10693 a_2162_n136236# a_2112_n66# a_1898_n136236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10694 a_2162_n127858# a_2112_n66# a_2030_n127858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10695 word304 A0 a_2294_n43368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10696 GND A8 word512 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10697 word713 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10698 a_1766_n37404# A3 a_1502_n37404# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10699 a_2294_n102014# A1 a_1898_n102014# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10700 word233 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10701 word976 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10702 a_1766_n132260# A3 a_1502_n132260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10703 word841 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10704 GND A2 word82 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10705 a_2030_n42658# A2 a_1634_n42658# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10706 a_578_n104854# a_528_n66# a_446_n104854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10707 GND A5 word513 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10708 GND A5 word454 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10709 GND A9 word506 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10710 a_2294_n49048# A1 a_2030_n49048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10711 a_710_n113516# A7 a_314_n113516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10712 a_1766_n109398# A3 a_1502_n109398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10713 word709 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10714 GND A9 word447 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10715 GND A4 word843 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10716 a_2162_n33570# a_2112_n66# a_2030_n33570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10717 GND A8 word27 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10718 word626 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10719 a_710_n37688# A7 a_314_n37688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10720 a_710_n46066# A7 a_314_n46066# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10721 word570 A0 a_2162_n81140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10722 a_2030_n19796# A2 a_1634_n19796# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10723 GND A8 word129 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10724 word754 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10725 a_1898_n118060# a_1848_n66# a_1634_n118060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10726 word628 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10727 a_1898_n140496# a_1848_n66# a_1634_n140496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10728 a_2294_n131408# A1 a_1898_n131408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10729 word777 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10730 a_446_n23346# A8 a_182_n23346# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10731 word499 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10732 a_1634_n97186# a_1584_n66# a_1502_n97186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10733 a_446_n14968# A8 a_182_n14968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10734 GND A1 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10735 GND A6 word58 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10736 word440 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10737 word350 A0 a_2162_n49900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10738 GND A8 word617 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10739 GND A9 word225 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10740 word759 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10741 GND A8 word746 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10742 GND A4 word779 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10743 a_578_n142626# a_528_n66# a_314_n142626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10744 a_446_n92642# A8 a_50_n92642# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10745 GND A6 word900 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10746 GND A6 word959 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10747 a_2294_n130982# A1 a_2030_n130982# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10748 GND A1 word820 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10749 GND A2 word187 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10750 a_446_n102440# A8 a_50_n102440# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10751 word765 a_2376_n66# a_2294_n108830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10752 a_2030_n126296# A2 a_1634_n126296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10753 a_578_n128142# a_528_n66# a_314_n128142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10754 a_1106_n4886# a_1056_n66# a_974_n4886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10755 a_710_n75460# A7 a_446_n75460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10756 word1020 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10757 word522 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10758 word645 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10759 a_2162_n142058# a_2112_n66# a_1898_n142058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10760 word729 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10761 word463 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10762 a_1766_n34848# A3 a_1370_n34848# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10763 GND A1 word329 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10764 GND A1 word876 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10765 GND A3 word821 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10766 word13 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10767 a_2162_n119196# a_2112_n66# a_1898_n119196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10768 word821 a_2376_n66# a_2294_n116782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10769 a_1106_n15820# a_1056_n66# a_842_n15820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10770 a_1370_n122462# a_1320_n66# a_1238_n122462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10771 word545 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10772 a_1502_n626# A4 a_1238_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10773 a_446_n29878# A8 a_182_n29878# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10774 word955 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10775 GND A9 word330 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10776 GND A4 word943 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10777 GND A5 word846 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10778 GND A5 word787 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10779 a_1106_n23772# a_1056_n66# a_974_n23772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10780 a_710_n110960# A7 a_314_n110960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10781 GND A8 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10782 GND A0 word924 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10783 GND A8 word170 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10784 a_1238_n129136# A5 a_974_n129136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10785 word238 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10786 word297 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10787 word227 a_2376_n66# a_2162_n32434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10788 word1011 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10789 GND A0 word146 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10790 word893 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10791 a_446_n20790# A8 a_182_n20790# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10792 GND A1 word104 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10793 GND A6 word40 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10794 word978 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10795 word450 A0 a_2162_n64100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10796 GND A8 word658 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10797 a_50_n119906# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10798 a_446_n76028# A8 a_50_n76028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10799 GND A8 word728 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10800 word859 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10801 GND A8 word226 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10802 a_2294_n114368# A1 a_1898_n114368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10803 word59 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10804 a_2162_n9572# a_2112_n66# a_2030_n9572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10805 a_1766_n80572# A3 a_1370_n80572# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10806 a_2294_n105990# A1 a_2030_n105990# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10807 GND A7 word28 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10808 a_1370_n79862# a_1320_n66# a_1106_n79862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10809 GND A8 word556 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10810 GND A3 word865 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10811 a_1106_n61544# a_1056_n66# a_974_n61544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10812 word789 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10813 a_1238_n120048# A5 a_842_n120048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10814 a_1238_n111670# A5 a_974_n111670# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10815 GND A4 word718 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10816 word865 a_2376_n66# a_2294_n123030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10817 GND A5 word600 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10818 word493 a_2376_n66# a_2294_n70206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10819 word504 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10820 GND A6 word681 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10821 GND A1 word429 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10822 GND A7 word289 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10823 a_1502_n137656# A4 a_1238_n137656# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10824 a_974_n3040# A6 a_710_n3040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10825 a_50_n110818# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10826 a_710_n125870# A7 a_314_n125870# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10827 a_1370_n48338# a_1320_n66# a_1238_n48338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10828 a_1370_n39960# a_1320_n66# a_1238_n39960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10829 a_1370_n70774# a_1320_n66# a_1106_n70774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10830 GND A7 word560 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10831 GND A0 word970 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10832 a_1766_n87530# A3 a_1502_n87530# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10833 word273 a_2376_n66# a_2294_n38966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10834 word923 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10835 word124 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10836 a_1766_n26186# A3 a_1370_n26186# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10837 GND A1 word209 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10838 GND A1 word268 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10839 a_446_n35700# A8 a_182_n35700# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10840 a_1106_n90938# a_1056_n66# a_842_n90938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10841 word962 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10842 GND A2 word435 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10843 GND A7 word616 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10844 a_2294_n129278# A1 a_1898_n129278# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10845 a_578_n21642# a_528_n66# a_446_n21642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10846 GND A5 word23 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10847 a_974_n60834# A6 a_578_n60834# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10848 word835 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10849 word894 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10850 GND A5 word726 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10851 a_578_n68502# a_528_n66# a_314_n68502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10852 a_1370_n86110# a_1320_n66# a_1238_n86110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10853 a_1502_n114084# A4 a_1106_n114084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10854 a_314_n41806# a_264_n66# a_182_n41806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10855 GND A1 word145 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10856 word668 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10857 a_1370_n16388# a_1320_n66# a_1106_n16388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10858 word539 a_2376_n66# a_2162_n76738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10859 GND A0 word804 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10860 a_446_n2330# A8 a_182_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10861 a_50_n125728# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10862 a_50_n134106# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10863 GND A7 word335 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10864 word107 a_2376_n66# a_2162_n15394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10865 a_842_n30872# a_792_n66# a_578_n30872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10866 a_974_n37972# A6 a_710_n37972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10867 a_1766_n55580# A3 a_1502_n55580# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10868 a_2294_n120190# A1 a_1898_n120190# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10869 a_1370_n94062# a_1320_n66# a_1238_n94062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10870 word756 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10871 a_182_n11844# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10872 a_182_n20222# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10873 a_1370_n85684# a_1320_n66# a_1238_n85684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10874 word236 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10875 GND A8 word538 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10876 word969 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10877 a_182_n58704# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10878 word446 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10879 a_50_n81708# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10880 word28 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10881 a_2294_n4318# A1 a_1898_n4318# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10882 GND A4 word229 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10883 a_1370_n54160# a_1320_n66# a_1106_n54160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10884 GND A5 word69 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10885 a_842_n46208# a_792_n66# a_710_n46208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10886 GND A0 word134 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10887 word373 a_2376_n66# a_2294_n53166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10888 a_974_n75744# A6 a_710_n75744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10889 a_182_n9004# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10890 a_50_n102156# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10891 GND A6 word561 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10892 word1022 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10893 a_314_n56716# a_264_n66# a_182_n56716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10894 GND A0 word292 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10895 GND A1 word309 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10896 word980 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10897 word1003 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10898 a_2030_n7016# A2 a_1766_n7016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10899 GND A0 word622 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10900 a_842_n45782# a_792_n66# a_710_n45782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10901 word948 A0 a_2294_n134816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10902 a_182_n35132# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10903 a_182_n26754# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10904 word221 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10905 a_974_n44220# A6 a_710_n44220# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10906 GND A6 word280 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10907 GND A0 word70 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10908 a_578_n65946# a_528_n66# a_314_n65946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10909 a_1898_n56432# a_1848_n66# a_1634_n56432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10910 word842 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10911 a_710_n7158# A7 a_446_n7158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10912 a_50_n96618# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10913 GND A3 word37 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10914 word47 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10915 word650 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10916 a_842_n14258# a_792_n66# a_710_n14258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10917 a_974_n111812# A6 a_710_n111812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10918 word831 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10919 a_50_n131550# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10920 word612 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10921 word772 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10922 a_1634_n33712# a_1584_n66# a_1502_n33712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10923 a_974_n43794# A6 a_710_n43794# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10924 GND A4 word393 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10925 word553 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10926 GND A4 word334 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10927 word424 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10928 a_974_n99032# A6 a_578_n99032# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10929 word738 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10930 GND A6 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10931 a_842_n83554# a_792_n66# a_710_n83554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10932 a_50_n117066# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10933 word419 a_2376_n66# a_2162_n59698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10934 word778 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10935 a_182_n64526# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10936 a_50_n108688# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10937 a_1502_n55012# A4 a_1238_n55012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10938 word782 A0 a_2162_n111244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10939 a_1502_n46634# A4 a_1238_n46634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10940 a_314_n117918# a_264_n66# a_50_n117918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10941 word263 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10942 GND A2 word640 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10943 a_1898_n94204# a_1848_n66# a_1766_n94204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10944 a_1502_n6306# A4 a_1106_n6306# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10945 word708 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10946 a_842_n122462# a_792_n66# a_710_n122462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10947 a_578_n33996# a_528_n66# a_446_n33996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10948 a_50_n73046# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10949 a_974_n59130# A6 a_578_n59130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10950 a_842_n52030# a_792_n66# a_710_n52030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10951 word324 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10952 a_974_n81566# A6 a_710_n81566# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10953 a_1106_n97186# a_1056_n66# a_974_n97186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10954 GND A6 word661 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10955 a_182_n6448# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10956 a_1502_n15110# A4 a_1106_n15110# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10957 a_314_n62538# a_264_n66# a_182_n62538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10958 word1004 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10959 GND A4 word109 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10960 GND A4 word168 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10961 GND A0 word950 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10962 a_1634_n112806# a_1584_n66# a_1370_n112806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10963 a_842_n29168# a_792_n66# a_578_n29168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10964 word685 a_2376_n66# a_2294_n97470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10965 GND A0 word604 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10966 a_314_n48054# a_264_n66# a_182_n48054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10967 word470 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10968 a_182_n32576# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10969 a_314_n39676# a_264_n66# a_182_n39676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10970 a_1502_n14684# A4 a_1106_n14684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10971 a_1502_n23062# A4 a_1106_n23062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10972 a_1106_n106132# a_1056_n66# a_842_n106132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10973 a_1370_n7016# a_1320_n66# a_1106_n7016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10974 a_578_n71768# a_528_n66# a_314_n71768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10975 a_1898_n62254# a_1848_n66# a_1766_n62254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10976 word883 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10977 GND A3 word279 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10978 word533 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10979 word592 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10980 word828 A0 a_2294_n117776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10981 GND A3 word496 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10982 a_182_n18092# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10983 GND A3 word19 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10984 word61 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10985 a_974_n27180# A6 a_578_n27180# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10986 word491 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10987 word872 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10988 GND A2 word944 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10989 word222 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10990 word813 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10991 a_578_n57284# a_528_n66# a_314_n57284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10992 a_1898_n39392# a_1848_n66# a_1766_n39392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X10993 a_1238_n47202# A5 a_842_n47202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10994 word594 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10995 a_842_n137372# a_792_n66# a_578_n137372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10996 a_1238_n38824# A5 a_974_n38824# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X10997 a_50_n79578# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10998 GND A4 word7 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X10999 a_974_n96476# A6 a_578_n96476# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11000 GND A0 word438 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11001 a_182_n70348# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11002 word201 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11003 GND A3 word215 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11004 a_1106_n135526# a_1056_n66# a_974_n135526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11005 a_182_n61970# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11006 a_314_n123740# a_264_n66# a_50_n123740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11007 a_314_n132118# a_264_n66# a_50_n132118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11008 word648 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11009 word304 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11010 word427 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11011 a_1898_n106842# a_1848_n66# a_1634_n106842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11012 GND A5 word212 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11013 a_1898_n91648# a_1848_n66# a_1766_n91648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11014 GND A5 word153 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11015 word157 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11016 GND A3 word113 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11017 word365 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11018 a_182_n47486# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11019 GND A2 word66 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11020 a_1502_n29594# A4 a_1238_n29594# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11021 a_314_n109256# a_264_n66# a_50_n109256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11022 word487 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11023 GND A9 word146 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11024 a_578_n95056# a_528_n66# a_446_n95056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11025 a_314_n131692# a_264_n66# a_50_n131692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11026 word266 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11027 a_1898_n77164# a_1848_n66# a_1634_n77164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11028 word697 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11029 word204 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11030 word327 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11031 a_974_n132544# A6 a_578_n132544# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11032 a_1634_n54444# a_1584_n66# a_1370_n54444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11033 word467 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11034 word699 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11035 GND A4 word480 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11036 a_2162_n108404# a_2112_n66# a_2030_n108404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11037 word108 A0 a_2294_n15536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11038 a_314_n45498# a_264_n66# a_182_n45498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11039 word692 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11040 a_1634_n104144# a_1584_n66# a_1370_n104144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11041 a_1370_n4460# a_1320_n66# a_1238_n4460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11042 word423 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11043 a_974_n109682# A6 a_710_n109682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11044 GND A3 word320 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11045 word596 A0 a_2294_n84832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11046 word633 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11047 word105 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11048 a_314_n138650# a_264_n66# a_50_n138650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11049 word591 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11050 word694 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11051 word409 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11052 word140 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11053 a_2030_n23204# A2 a_1766_n23204# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11054 word350 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11055 GND A2 word985 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11056 word854 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11057 GND A5 word258 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11058 word635 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11059 a_842_n143194# a_792_n66# a_578_n143194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11060 word593 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11061 GND A7 word841 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11062 a_50_n85400# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11063 a_2162_n14116# a_2112_n66# a_2030_n14116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11064 GND A9 word251 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11065 a_1634_n83838# a_1584_n66# a_1502_n83838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11066 a_1634_n92216# a_1584_n66# a_1502_n92216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11067 a_710_n18234# A7 a_446_n18234# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11068 word102 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11069 word374 A0 a_2162_n53308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11070 a_1634_n22494# a_1584_n66# a_1370_n22494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11071 a_1106_n141348# a_1056_n66# a_842_n141348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11072 word7 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11073 word310 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11074 a_2162_n83412# a_2112_n66# a_2030_n83412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11075 a_1634_n133538# a_1584_n66# a_1502_n133538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11076 a_1106_n132970# a_1056_n66# a_974_n132970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11077 word716 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11078 word303 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11079 GND A6 word924 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11080 word244 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11081 a_1502_n96760# A4 a_1106_n96760# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11082 GND A7 word777 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11083 a_2294_n12128# A1 a_1898_n12128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11084 a_314_n115078# a_264_n66# a_50_n115078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11085 a_2030_n112948# A2 a_1634_n112948# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11086 word366 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11087 GND A5 word524 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11088 word469 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11089 word307 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11090 a_578_n92500# a_528_n66# a_446_n92500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11091 a_1238_n82418# A5 a_842_n82418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11092 GND A5 word92 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11093 GND A3 word642 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11094 a_1766_n119338# A3 a_1502_n119338# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11095 a_1238_n21074# A5 a_974_n21074# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11096 a_2294_n81424# A1 a_1898_n81424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11097 GND A3 word583 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11098 GND A6 word921 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11099 a_1238_n12696# A5 a_842_n12696# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11100 a_710_n47628# A7 a_314_n47628# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11101 a_2030_n38114# A2 a_1634_n38114# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11102 word368 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11103 a_1766_n141774# A3 a_1502_n141774# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11104 GND A3 word786 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11105 a_2030_n29736# A2 a_1766_n29736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11106 word959 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11107 word900 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11108 a_1634_n51888# a_1584_n66# a_1502_n51888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11109 word449 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11110 word765 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11111 a_2162_n114226# a_2112_n66# a_2030_n114226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11112 word90 A0 a_2162_n12980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11113 a_2162_n29026# a_2112_n66# a_2030_n29026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11114 a_1238_n81992# A5 a_842_n81992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11115 a_1634_n101588# a_1584_n66# a_1502_n101588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11116 a_446_n24908# A8 a_182_n24908# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11117 word510 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11118 word347 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11119 word207 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11120 word415 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11121 word420 A0 a_2294_n59840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11122 a_1502_n73188# A4 a_1238_n73188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11123 word829 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11124 a_2162_n98322# a_2112_n66# a_2030_n98322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11125 word450 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11126 a_1766_n110250# A3 a_1502_n110250# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11127 a_2030_n20648# A2 a_1766_n20648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11128 word566 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11129 GND A7 word882 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11130 a_842_n9856# a_792_n66# a_710_n9856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11131 word634 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11132 GND A9 word351 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11133 GND A9 word134 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11134 a_2294_n27038# A1 a_1898_n27038# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11135 a_2030_n67508# A2 a_1634_n67508# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11136 word476 A0 a_2294_n67792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11137 GND A9 word292 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11138 a_2030_n127858# A2 a_1766_n127858# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11139 a_578_n129704# a_528_n66# a_314_n129704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11140 word471 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11141 a_2162_n143620# a_2112_n66# a_2030_n143620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11142 a_710_n15678# A7 a_446_n15678# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11143 GND A5 word197 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11144 word943 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11145 GND A5 word138 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11146 word283 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11147 a_2162_n58420# a_2112_n66# a_2030_n58420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11148 a_2294_n96334# A1 a_1898_n96334# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11149 GND A3 word688 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11150 a_2162_n4602# a_2112_n66# a_1898_n4602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11151 word473 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11152 word613 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11153 word891 a_2376_n66# a_2162_n126722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11154 a_710_n84974# A7 a_446_n84974# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11155 word254 A0 a_2162_n36268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11156 GND A9 word70 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11157 word190 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11158 a_2162_n57994# a_2112_n66# a_1898_n57994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11159 a_2162_n66372# a_2112_n66# a_2030_n66372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11160 word615 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11161 a_974_n6732# A6 a_710_n6732# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11162 word183 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11163 a_1502_n88098# A4 a_1106_n88098# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11164 GND A1 word724 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11165 GND A6 word804 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11166 a_1766_n125160# A3 a_1370_n125160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11167 GND A2 word91 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11168 a_1106_n33712# a_1056_n66# a_842_n33712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11169 a_710_n53450# A7 a_314_n53450# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11170 a_578_n106132# a_528_n66# a_446_n106132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11171 word678 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11172 a_2030_n35558# A2 a_1634_n35558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11173 GND A5 word404 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11174 word865 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11175 word1000 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11176 word367 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11177 a_1238_n65378# A5 a_842_n65378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11178 a_1238_n57000# A5 a_974_n57000# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11179 word718 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11180 GND A7 word93 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11181 a_1502_n109824# A4 a_1238_n109824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11182 GND A9 word397 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11183 a_446_n30730# A8 a_182_n30730# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11184 a_1766_n21216# A3 a_1370_n21216# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11185 a_2294_n64384# A1 a_1898_n64384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11186 GND A1 word721 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11187 word520 A0 a_2294_n74040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11188 GND A9 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11189 word206 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11190 word929 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11191 GND A8 word237 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11192 GND A7 word581 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11193 a_446_n16246# A8 a_182_n16246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11194 a_1370_n89802# a_1320_n66# a_1106_n89802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11195 GND A7 word39 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11196 GND A9 word175 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11197 GND A2 word298 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11198 GND A7 word864 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11199 a_1238_n121610# A5 a_842_n121610# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11200 a_2030_n73330# A2 a_1766_n73330# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11201 a_1502_n100736# A4 a_1238_n100736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11202 a_1370_n138934# a_1320_n66# a_1238_n138934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11203 a_578_n135526# a_528_n66# a_314_n135526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11204 a_446_n85542# A8 a_50_n85542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11205 GND A5 word670 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11206 word574 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11207 GND A6 word909 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11208 GND A5 word962 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11209 word925 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11210 word142 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11211 GND A3 word932 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11212 a_1106_n6164# a_1056_n66# a_974_n6164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11213 GND A2 word137 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11214 a_1766_n50610# A3 a_1502_n50610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11215 word856 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11216 GND A1 word928 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11217 word472 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11218 a_2030_n81282# A2 a_1634_n81282# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11219 word595 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11220 word413 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11221 a_710_n90796# A7 a_446_n90796# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11222 a_1370_n80714# a_1320_n66# a_1106_n80714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11223 a_1370_n107410# a_1320_n66# a_1106_n107410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11224 GND A8 word562 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11225 a_2162_n126580# a_2112_n66# a_2030_n126580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11226 word343 a_2376_n66# a_2162_n48906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11227 word764 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11228 GND A8 word71 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11229 a_2294_n79294# A1 a_1898_n79294# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11230 a_1766_n27748# A3 a_1502_n27748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11231 GND A1 word496 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11232 a_2162_n72194# a_2112_n66# a_2030_n72194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11233 GND A7 word356 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11234 a_446_n103292# A8 a_50_n103292# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11235 GND A3 word771 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11236 GND A9 word54 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11237 word771 a_2376_n66# a_2162_n109682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11238 a_1370_n57852# a_1320_n66# a_1238_n57852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11239 GND A2 word505 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11240 GND A3 word710 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11241 word975 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11242 GND A2 word73 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11243 a_578_n103576# a_528_n66# a_446_n103576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11244 a_1370_n106984# a_1320_n66# a_1106_n106984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11245 a_2030_n41380# A2 a_1766_n41380# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11246 word905 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11247 a_1238_n136520# A5 a_842_n136520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11248 GND A5 word796 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11249 GND A2 word403 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11250 a_1502_n124024# A4 a_1106_n124024# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11251 GND A4 word834 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11252 GND A7 word75 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11253 a_710_n112238# A7 a_314_n112238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11254 GND A9 word438 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11255 a_1502_n115646# A4 a_1106_n115646# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11256 a_1106_n16672# a_1056_n66# a_842_n16672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11257 GND A3 word707 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11258 a_1370_n26328# a_1320_n66# a_1106_n26328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11259 word707 a_2376_n66# a_2162_n100594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11260 a_2294_n138792# A1 a_2030_n138792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11261 GND A0 word874 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11262 a_1370_n17950# a_1320_n66# a_1106_n17950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11263 GND A8 word120 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11264 word177 a_2376_n66# a_2294_n25334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11265 word188 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11266 word619 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11267 word961 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11268 a_446_n22068# A8 a_182_n22068# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11269 GND A0 word96 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11270 GND A1 word113 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11271 GND A6 word49 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11272 a_446_n13690# A8 a_182_n13690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11273 GND A8 word608 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11274 word809 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11275 GND A8 word176 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11276 a_1370_n144756# a_1320_n66# a_1106_n144756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11277 a_578_n141348# a_528_n66# a_314_n141348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11278 a_578_n132970# a_528_n66# a_314_n132970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11279 a_1766_n73472# A3 a_1502_n73472# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11280 a_446_n91364# A8 a_50_n91364# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11281 GND A1 word601 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11282 a_446_n82986# A8 a_50_n82986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11283 GND A6 word950 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11284 GND A2 word610 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11285 a_1106_n54444# a_1056_n66# a_842_n54444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11286 a_1238_n104570# A5 a_842_n104570# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11287 GND A2 word178 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11288 GND A6 word301 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11289 a_2030_n56290# A2 a_1634_n56290# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11290 a_710_n1762# A7 a_446_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11291 word443 a_2376_n66# a_2162_n63106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11292 GND A5 word901 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11293 word720 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11294 GND A5 word842 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11295 a_710_n127148# A7 a_314_n127148# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11296 a_50_n103718# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11297 GND A0 word362 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11298 GND A2 word666 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11299 a_710_n118770# A7 a_314_n118770# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11300 GND A1 word320 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11301 GND A8 word64 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11302 a_1370_n72052# a_1320_n66# a_1106_n72052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11303 a_1370_n63674# a_1320_n66# a_1106_n63674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11304 a_2294_n145040# A1 a_1898_n145040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11305 word873 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11306 a_1370_n121184# a_1320_n66# a_1238_n121184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11307 word814 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11308 a_446_n28600# A8 a_182_n28600# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11309 a_1502_n18802# A4 a_1238_n18802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11310 a_1766_n19086# A3 a_1502_n19086# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11311 GND A1 word45 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11312 GND A1 word376 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11313 GND A6 word567 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11314 GND A0 word976 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11315 GND A4 word875 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11316 GND A5 word778 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11317 GND A2 word385 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11318 a_710_n8720# A7 a_446_n8720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11319 GND A4 word74 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11320 a_446_n97896# A8 a_50_n97896# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11321 a_842_n15820# a_792_n66# a_710_n15820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11322 a_974_n62112# A6 a_578_n62112# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11323 word286 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11324 a_1106_n69354# a_1056_n66# a_842_n69354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11325 a_1238_n119480# A5 a_842_n119480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11326 word159 a_2376_n66# a_2162_n22778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11327 GND A6 word406 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11328 word1002 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11329 word867 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11330 word1019 a_2376_n66# a_2162_n144898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11331 word808 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11332 word825 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11333 GND A4 word36 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11334 word559 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11335 GND A0 word754 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11336 GND A8 word649 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11337 a_50_n127006# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11338 word489 a_2376_n66# a_2294_n69638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11339 GND A7 word344 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11340 GND A8 word590 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11341 a_50_n118628# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11342 GND A8 word719 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11343 a_1766_n48480# A3 a_1370_n48480# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11344 word498 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11345 a_182_n13122# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11346 a_974_n22210# A6 a_578_n22210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11347 GND A6 word184 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11348 a_1106_n60266# a_1056_n66# a_974_n60266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11349 word186 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11350 word746 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11351 a_1370_n136094# a_1320_n66# a_1106_n136094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11352 GND A2 word219 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11353 a_1106_n51888# a_1056_n66# a_842_n51888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11354 a_446_n3182# A8 a_182_n3182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11355 a_50_n74608# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11356 a_1898_n8862# a_1848_n66# a_1634_n8862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11357 word495 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11358 a_974_n91506# A6 a_578_n91506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11359 word425 a_2376_n66# a_2294_n60550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11360 GND A2 word490 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11361 a_1106_n98748# a_1056_n66# a_974_n98748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11362 GND A6 word672 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11363 a_1502_n128000# A4 a_1238_n128000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11364 a_578_n29452# a_528_n66# a_446_n29452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11365 a_974_n21784# A6 a_578_n21784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11366 word4 A0 a_2294_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11367 word41 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11368 GND A0 word1020 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11369 a_974_n77022# A6 a_710_n77022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11370 word323 a_2376_n66# a_2162_n46066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11371 word391 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11372 GND A0 word674 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11373 word115 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11374 GND A0 word242 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11375 GND A7 word119 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11376 a_182_n42516# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11377 a_314_n49616# a_264_n66# a_182_n49616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11378 a_1502_n24624# A4 a_1106_n24624# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11379 GND A1 word200 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11380 a_1502_n33002# A4 a_1106_n33002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11381 GND A8 word695 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11382 word603 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11383 word662 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11384 GND A7 word607 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11385 word898 A0 a_2162_n127716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11386 word806 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11387 a_578_n20364# a_528_n66# a_446_n20364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11388 a_1766_n9572# A3 a_1502_n9572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11389 a_842_n100452# a_792_n66# a_578_n100452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11390 GND A1 word688 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11391 a_182_n28032# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11392 a_974_n768# A6 a_710_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11393 a_974_n37120# A6 a_710_n37120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11394 a_182_n19654# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11395 word15 a_2376_n66# a_2162_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11396 GND A5 word14 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11397 word110 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11398 a_842_n30020# a_792_n66# a_578_n30020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11399 GND A2 word955 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11400 a_578_n67224# a_528_n66# a_314_n67224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11401 a_578_n58846# a_528_n66# a_314_n58846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11402 GND A6 word447 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11403 a_842_n138934# a_792_n66# a_578_n138934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11404 a_314_n40528# a_264_n66# a_182_n40528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11405 a_50_n89518# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11406 word56 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11407 word600 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11408 a_842_n90938# a_792_n66# a_710_n90938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11409 a_50_n124450# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11410 word166 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11411 a_1634_n26612# a_1584_n66# a_1370_n26612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11412 a_974_n36694# A6 a_710_n36694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11413 a_974_n45072# A6 a_710_n45072# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11414 GND A0 word508 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11415 GND A2 word1011 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11416 a_182_n71910# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11417 word747 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11418 word374 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11419 word315 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11420 a_182_n10566# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11421 word227 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11422 a_842_n107410# a_792_n66# a_578_n107410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11423 a_1898_n31866# a_1848_n66# a_1634_n31866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11424 a_182_n57426# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11425 a_50_n80430# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11426 word378 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11427 word437 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11428 GND A6 word555 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11429 word732 A0 a_2294_n104144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11430 a_2294_n3040# A1 a_1898_n3040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11431 a_578_n96618# a_528_n66# a_446_n96618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11432 a_314_n141632# a_264_n66# a_50_n141632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11433 a_1898_n87104# a_1848_n66# a_1766_n87104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11434 word717 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11435 word371 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11436 a_1502_n142200# A4 a_1106_n142200# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11437 GND A2 word730 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11438 word911 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11439 a_578_n35274# a_528_n66# a_446_n35274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11440 a_578_n26896# a_528_n66# a_446_n26896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11441 word276 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11442 a_842_n106984# a_792_n66# a_578_n106984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11443 a_974_n74466# A6 a_710_n74466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11444 GND A6 word552 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11445 word954 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11446 word1013 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11447 a_314_n55438# a_264_n66# a_182_n55438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11448 a_314_n110108# a_264_n66# a_50_n110108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11449 word493 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11450 a_50_n139360# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11451 word434 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11452 word994 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11453 word271 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11454 GND A0 word554 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11455 word935 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11456 word847 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11457 a_1502_n68928# A4 a_1106_n68928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11458 word479 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11459 GND A4 word547 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11460 word420 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11461 a_182_n25476# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11462 word924 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11463 word111 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11464 a_578_n64668# a_528_n66# a_314_n64668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11465 word542 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11466 a_842_n144756# a_792_n66# a_578_n144756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11467 a_50_n95340# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11468 word38 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11469 word231 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11470 word639 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11471 a_974_n110534# A6 a_710_n110534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11472 word476 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11473 GND A2 word835 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11474 a_1766_n113942# A3 a_1502_n113942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11475 word544 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11476 word763 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11477 GND A4 word325 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11478 word921 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11479 a_1106_n142910# a_1056_n66# a_842_n142910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11480 word18 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11481 a_1898_n122604# a_1848_n66# a_1634_n122604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11482 a_842_n82276# a_792_n66# a_710_n82276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11483 GND A3 word224 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11484 GND A0 word388 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11485 a_182_n54870# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11486 a_182_n63248# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11487 GND A3 word165 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11488 a_314_n125018# a_264_n66# a_50_n125018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11489 word714 A0 a_2162_n101588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11490 word6 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11491 a_1502_n36978# A4 a_1238_n36978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11492 a_314_n116640# a_264_n66# a_50_n116640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11493 a_1502_n5028# A4 a_1106_n5028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11494 a_710_n10708# A7 a_446_n10708# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11495 a_1238_n31014# A5 a_842_n31014# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11496 a_842_n121184# a_792_n66# a_710_n121184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11497 a_1238_n22636# A5 a_974_n22636# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11498 a_2030_n108404# A2 a_1634_n108404# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11499 a_1634_n70206# a_1584_n66# a_1502_n70206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11500 a_974_n80288# A6 a_710_n80288# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11501 word970 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11502 GND A9 word96 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11503 a_314_n124592# a_264_n66# a_50_n124592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11504 a_182_n5170# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11505 word995 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11506 a_314_n61260# a_264_n66# a_182_n61260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11507 word87 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11508 word160 A0 a_2294_n22920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11509 GND A3 word551 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11510 a_1238_n91932# A5 a_974_n91932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11511 GND A4 word100 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11512 word155 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11513 a_2162_n61402# a_2112_n66# a_1898_n61402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11514 a_2294_n68502# A1 a_2030_n68502# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11515 GND A0 word654 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11516 a_1634_n47344# a_1584_n66# a_1502_n47344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11517 word417 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11518 a_1502_n83128# A4 a_1238_n83128# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11519 word55 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11520 a_1502_n74750# A4 a_1238_n74750# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11521 word891 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11522 a_314_n38398# a_264_n66# a_182_n38398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11523 GND A4 word588 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11524 word643 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11525 GND A4 word647 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11526 a_1898_n137514# a_1848_n66# a_1766_n137514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11527 a_182_n31298# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11528 word216 A0 a_2294_n30872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11529 word211 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11530 word636 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11531 a_578_n70490# a_528_n66# a_314_n70490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11532 a_182_n69780# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11533 word546 A0 a_2162_n77732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11534 GND A9 word362 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11535 GND A0 word42 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11536 word52 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11537 a_2030_n16104# A2 a_1766_n16104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11538 word213 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11539 word482 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11540 word804 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11541 GND A5 word208 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11542 GND A5 word267 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11543 word353 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11544 word585 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11545 word745 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11546 a_1238_n37546# A5 a_974_n37546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11547 a_50_n78300# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11548 GND A3 word326 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11549 a_974_n95198# A6 a_578_n95198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11550 word484 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11551 GND A9 word201 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11552 a_2294_n36552# A1 a_2030_n36552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11553 word355 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11554 word519 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11555 a_1634_n76738# a_1584_n66# a_1370_n76738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11556 word324 A0 a_2294_n46208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11557 a_1634_n15394# a_1584_n66# a_1502_n15394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11558 a_1502_n51178# A4 a_1106_n51178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11559 a_1106_n134248# a_1056_n66# a_974_n134248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11560 a_1634_n126438# a_1584_n66# a_1370_n126438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11561 a_1502_n42800# A4 a_1106_n42800# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11562 word295 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11563 a_1106_n125870# a_1056_n66# a_842_n125870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11564 a_1898_n105564# a_1848_n66# a_1766_n105564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11565 word253 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11566 GND A0 word700 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11567 GND A5 word144 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11568 GND A6 word815 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11569 a_2030_n114226# A2 a_1766_n114226# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11570 GND A2 word57 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11571 GND A5 word474 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11572 a_2030_n105848# A2 a_1634_n105848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11573 word478 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11574 word419 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11575 a_2162_n121610# a_2112_n66# a_1898_n121610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11576 a_1238_n66940# A5 a_842_n66940# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11577 a_1238_n75318# A5 a_974_n75318# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11578 word729 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11579 a_2162_n36410# a_2112_n66# a_1898_n36410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11580 GND A3 word592 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11581 GND A9 word467 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11582 GND A3 word533 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11583 GND A3 word736 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11584 a_1766_n134674# A3 a_1370_n134674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11585 word909 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11586 a_974_n131266# A6 a_578_n131266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11587 a_1634_n44788# a_1584_n66# a_1370_n44788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11588 word399 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11589 word690 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11590 a_1238_n74892# A5 a_974_n74892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11591 a_1898_n134958# a_1848_n66# a_1766_n134958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11592 a_446_n17808# A8 a_182_n17808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11593 a_2162_n44362# a_2112_n66# a_1898_n44362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11594 a_1766_n103150# A3 a_1370_n103150# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11595 a_2030_n143620# A2 a_1766_n143620# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11596 word523 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11597 word685 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11598 word845 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11599 a_2294_n133822# A1 a_1898_n133822# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11600 word710 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11601 word153 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11602 GND A7 word832 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11603 word584 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11604 GND A7 word773 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11605 a_1106_n7726# a_1056_n66# a_974_n7726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11606 a_2030_n91222# A2 a_1766_n91222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11607 word665 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11608 GND A9 word242 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11609 a_2294_n42374# A1 a_2030_n42374# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11610 word233 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11611 a_1370_n20932# a_1320_n66# a_1238_n20932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11612 word715 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11613 GND A8 word82 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11614 GND A8 word141 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11615 a_2162_n73756# a_2112_n66# a_1898_n73756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11616 GND A1 word896 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11617 word707 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11618 a_1634_n68076# a_1584_n66# a_1370_n68076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11619 a_446_n104854# A8 a_50_n104854# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11620 word841 a_2376_n66# a_2294_n119622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11621 a_1898_n111386# a_1848_n66# a_1634_n111386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11622 word235 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11623 a_710_n77874# A7 a_446_n77874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11624 a_710_n86252# A7 a_446_n86252# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11625 GND A6 word915 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11626 word204 A0 a_2294_n29168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11627 GND A6 word11 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11628 a_1370_n125302# a_1320_n66# a_1106_n125302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11629 word843 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11630 a_1370_n116924# a_1320_n66# a_1106_n116924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11631 a_2030_n51320# A2 a_1634_n51320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11632 GND A5 word515 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11633 a_2030_n111670# A2 a_1766_n111670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11634 a_2294_n101872# A1 a_1898_n101872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11635 word692 A0 a_2294_n98464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11636 GND A9 word508 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11637 GND A9 word449 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11638 a_1106_n26612# a_1056_n66# a_974_n26612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11639 GND A8 word29 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11640 a_710_n46350# A7 a_314_n46350# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11641 word499 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11642 a_2294_n71768# A1 a_2030_n71768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11643 word359 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11644 word950 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11645 word317 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11646 word621 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11647 word777 a_2376_n66# a_2294_n110534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11648 a_1238_n58278# A5 a_974_n58278# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11649 a_2162_n104570# a_2112_n66# a_1898_n104570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11650 word140 A0 a_2294_n20080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11651 a_1238_n49900# A5 a_842_n49900# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11652 word630 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11653 GND A9 word347 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11654 word779 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11655 a_446_n32008# A8 a_182_n32008# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11656 a_1766_n14116# A3 a_1502_n14116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11657 a_2162_n19370# a_2112_n66# a_1898_n19370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11658 a_1634_n97470# a_1584_n66# a_1502_n97470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11659 a_1898_n140780# a_1848_n66# a_1634_n140780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11660 a_446_n23630# A8 a_182_n23630# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11661 GND A6 word60 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11662 GND A1 word124 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11663 a_710_n121752# A7 a_314_n121752# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11664 GND A8 word26 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11665 word1012 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11666 word879 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11667 a_1370_n35842# a_1320_n66# a_1106_n35842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11668 GND A8 word246 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11669 GND A7 word531 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11670 GND A8 word748 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11671 a_578_n142910# a_528_n66# a_314_n142910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11672 GND A8 word187 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11673 a_2162_n88666# a_2112_n66# a_1898_n88666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11674 a_2162_n97044# a_2112_n66# a_2030_n97044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11675 a_2294_n117208# A1 a_2030_n117208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11676 a_446_n92926# A8 a_50_n92926# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11677 a_2294_n108830# A1 a_1898_n108830# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11678 GND A7 word48 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11679 a_446_n31582# A8 a_182_n31582# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11680 GND A7 word873 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11681 GND A2 word248 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11682 a_2030_n66230# A2 a_1766_n66230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11683 a_1502_n102014# A4 a_1238_n102014# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11684 GND A7 word814 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11685 GND A9 word283 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11686 a_2030_n126580# A2 a_1634_n126580# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11687 a_578_n128426# a_528_n66# a_314_n128426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11688 a_446_n78442# A8 a_50_n78442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11689 word524 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11690 a_710_n14400# A7 a_446_n14400# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11691 GND A5 word912 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11692 a_2294_n116782# A1 a_1898_n116782# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11693 word92 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11694 a_974_n25902# A6 a_578_n25902# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11695 a_1766_n43510# A3 a_1370_n43510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11696 a_2294_n86678# A1 a_2030_n86678# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11697 word464 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11698 a_2294_n95056# A1 a_1898_n95056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11699 word806 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11700 GND A1 word937 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11701 GND A3 word882 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11702 a_1238_n122462# A5 a_842_n122462# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11703 word15 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11704 a_2162_n3324# a_2112_n66# a_1898_n3324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11705 a_710_n83696# A7 a_446_n83696# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11706 a_2030_n74182# A2 a_1634_n74182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11707 word545 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11708 word1019 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11709 word943 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11710 a_1370_n131124# a_1320_n66# a_1238_n131124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11711 a_1370_n122746# a_1320_n66# a_1238_n122746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11712 word787 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11713 GND A7 word306 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11714 GND A0 word716 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11715 a_1502_n910# A4 a_1238_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11716 a_974_n5454# A6 a_710_n5454# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11717 GND A9 word63 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11718 GND A5 word848 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11719 GND A6 word795 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11720 a_1106_n32434# a_1056_n66# a_842_n32434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11721 a_1766_n98322# A3 a_1370_n98322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11722 a_1370_n108262# a_1320_n66# a_1106_n108262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11723 a_2030_n34280# A2 a_1766_n34280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11724 GND A6 word146 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11725 GND A5 word395 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11726 word299 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11727 a_1238_n64100# A5 a_842_n64100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11728 a_1238_n129420# A5 a_974_n129420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11729 word229 a_2376_n66# a_2294_n32718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11730 GND A7 word84 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11731 GND A9 word388 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11732 GND A1 word165 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11733 GND A1 word224 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11734 GND A4 word1001 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11735 GND A4 word942 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11736 a_1766_n11560# A3 a_1370_n11560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11737 GND A0 word824 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11738 a_1370_n50042# a_1320_n66# a_1238_n50042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11739 word980 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11740 GND A8 word660 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11741 word138 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11742 GND A7 word572 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11743 word127 a_2376_n66# a_2162_n18234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11744 a_842_n33712# a_792_n66# a_578_n33712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11745 GND A8 word228 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11746 word718 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11747 GND A8 word730 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11748 word911 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11749 a_1238_n137372# A5 a_842_n137372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11750 a_2294_n123030# A1 a_2030_n123030# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11751 a_2030_n89092# A2 a_1766_n89092# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11752 GND A1 word653 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11753 a_1238_n128994# A5 a_974_n128994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11754 GND A1 word221 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11755 GND A7 word30 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11756 a_1106_n70206# a_1056_n66# a_842_n70206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11757 GND A8 word558 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11758 word951 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11759 word892 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11760 GND A2 word289 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11761 a_1106_n61828# a_1056_n66# a_974_n61828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11762 a_578_n134248# a_528_n66# a_314_n134248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11763 word14 A0 a_2162_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11764 GND A8 word126 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11765 a_446_n4744# A8 a_182_n4744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11766 word48 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11767 a_446_n75886# A8 a_50_n75886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11768 a_446_n84264# A8 a_50_n84264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11769 a_1766_n66372# A3 a_1370_n66372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11770 a_1766_n57994# A3 a_1370_n57994# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11771 GND A2 word560 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11772 a_974_n40102# A6 a_710_n40102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11773 a_1502_n137940# A4 a_1238_n137940# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11774 GND A2 word128 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11775 word847 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11776 a_2030_n49190# A2 a_1634_n49190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11777 word923 a_2376_n66# a_2162_n131266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11778 GND A3 word864 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11779 GND A4 word776 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11780 word393 a_2376_n66# a_2294_n56006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11781 word925 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11782 GND A0 word312 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11783 GND A2 word616 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11784 a_974_n2898# A6 a_710_n2898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11785 GND A1 word428 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11786 GND A9 word45 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11787 a_842_n48622# a_792_n66# a_710_n48622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11788 word726 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11789 GND A7 word618 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11790 word764 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11791 a_578_n21926# a_528_n66# a_446_n21926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11792 a_578_n30304# a_528_n66# a_446_n30304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11793 a_1898_n12412# a_1848_n66# a_1766_n12412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11794 word241 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11795 a_578_n102298# a_528_n66# a_446_n102298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11796 a_1766_n95766# A3 a_1502_n95766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11797 GND A5 word25 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11798 GND A5 word728 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11799 GND A2 word394 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11800 GND A6 word517 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11801 a_1502_n114368# A4 a_1106_n114368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11802 a_1106_n15394# a_1056_n66# a_842_n15394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11803 a_446_n99174# A8 a_50_n99174# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11804 a_1502_n105990# A4 a_1106_n105990# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11805 word670 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11806 word236 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11807 a_974_n55012# A6 a_578_n55012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11808 word109 a_2376_n66# a_2294_n15678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11809 word952 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11810 word969 a_2376_n66# a_2294_n137798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11811 word817 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11812 word758 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11813 a_182_n20506# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11814 a_710_n9572# A7 a_446_n9572# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11815 GND A4 word512 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11816 a_1370_n85968# a_1320_n66# a_1238_n85968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11817 a_1370_n94346# a_1320_n66# a_1238_n94346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11818 GND A8 word599 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11819 GND A8 word540 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11820 a_1370_n143478# a_1320_n66# a_1106_n143478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11821 word798 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11822 a_578_n140070# a_528_n66# a_314_n140070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11823 a_842_n16672# a_792_n66# a_710_n16672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11824 a_50_n142342# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11825 a_1898_n41806# a_1848_n66# a_1766_n41806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11826 word597 a_2376_n66# a_2294_n84974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11827 a_50_n133964# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11828 word30 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11829 a_446_n90086# A8 a_50_n90086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11830 GND A1 word533 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11831 GND A1 word592 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11832 GND A6 word134 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11833 word136 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11834 word441 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11835 word981 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11836 GND A2 word169 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11837 a_1898_n27322# a_1848_n66# a_1634_n27322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11838 a_1106_n44788# a_1056_n66# a_974_n44788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11839 a_1106_n53166# a_1056_n66# a_842_n53166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11840 a_842_n125302# a_792_n66# a_710_n125302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11841 a_1898_n18944# a_1848_n66# a_1766_n18944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11842 GND A6 word292 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11843 word346 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11844 word445 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11845 GND A5 word833 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11846 a_974_n23062# A6 a_578_n23062# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11847 word375 a_2376_n66# a_2162_n53450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11848 a_1502_n129278# A4 a_1238_n129278# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11849 a_50_n102440# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11850 GND A0 word294 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11851 GND A2 word657 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11852 GND A2 word856 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11853 GND A4 word129 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11854 a_842_n54444# a_792_n66# a_710_n54444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11855 word341 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11856 a_1370_n62396# a_1320_n66# a_1106_n62396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11857 GND A0 word624 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11858 word917 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11859 a_1898_n1052# a_1848_n66# a_1766_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11860 GND A0 word192 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11861 word282 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11862 GND A4 word617 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11863 a_182_n8862# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11864 a_182_n35416# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11865 a_50_n110392# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11866 word223 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11867 a_314_n64952# a_264_n66# a_182_n64952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11868 word903 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11869 a_1898_n56716# a_1848_n66# a_1634_n56716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11870 GND A7 word557 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11871 a_1502_n120190# A4 a_1238_n120190# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11872 GND A1 word697 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11873 word756 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11874 GND A3 word39 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11875 word121 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11876 GND A2 word905 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11877 a_1106_n59698# a_1056_n66# a_974_n59698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11878 GND A6 word397 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11879 word991 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11880 a_974_n99316# A6 a_578_n99316# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11881 GND A6 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11882 a_842_n83838# a_792_n66# a_710_n83838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11883 GND A8 word640 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11884 a_50_n117350# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11885 a_1898_n8010# a_1848_n66# a_1766_n8010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11886 GND A0 word458 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11887 word21 a_2376_n66# a_2294_n3182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11888 word116 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11889 a_1634_n19512# a_1584_n66# a_1502_n19512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11890 GND A2 word961 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11891 word784 A0 a_2294_n111528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11892 a_182_n64810# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11893 a_1502_n46918# A4 a_1238_n46918# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11894 GND A1 word633 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11895 word611 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11896 word324 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11897 GND A4 word392 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11898 GND A4 word451 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11899 word265 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11900 GND A6 word175 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11901 a_842_n69354# a_792_n66# a_578_n69354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11902 word177 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11903 word1022 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11904 a_1898_n7584# a_1848_n66# a_1766_n7584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11905 a_1898_n24766# a_1848_n66# a_1634_n24766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11906 a_842_n122746# a_792_n66# a_710_n122746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11907 a_50_n73330# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11908 GND A3 word291 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11909 a_182_n72762# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11910 a_974_n81850# A6 a_710_n81850# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11911 a_314_n134532# a_264_n66# a_50_n134532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11912 a_1106_n97470# a_1056_n66# a_974_n97470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11913 GND A6 word663 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11914 GND A2 word739 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11915 word321 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11916 a_1634_n10424# a_1584_n66# a_1502_n10424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11917 a_842_n108262# a_792_n66# a_578_n108262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11918 a_578_n19796# a_528_n66# a_446_n19796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11919 a_578_n28174# a_528_n66# a_446_n28174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11920 GND A4 word170 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11921 a_50_n81282# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11922 word382 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11923 a_842_n51888# a_792_n66# a_710_n51888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11924 a_974_n58988# A6 a_578_n58988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11925 a_182_n32860# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11926 a_314_n39960# a_264_n66# a_182_n39960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11927 a_182_n41238# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11928 a_314_n48338# a_264_n66# a_182_n48338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11929 a_1502_n23346# A4 a_1106_n23346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11930 word286 A0 a_2162_n40812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11931 a_1106_n106416# a_1056_n66# a_842_n106416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11932 word443 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11933 a_314_n70774# a_264_n66# a_182_n70774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11934 a_1502_n14968# A4 a_1106_n14968# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11935 GND A4 word226 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11936 word384 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11937 word222 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11938 a_1898_n62538# a_1848_n66# a_1766_n62538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11939 a_1238_n1052# A5 a_974_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11940 word594 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11941 word797 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11942 GND A3 word498 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11943 GND A4 word556 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11944 a_1502_n92642# A4 a_1238_n92642# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11945 a_182_n18376# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11946 word874 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11947 word815 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11948 word655 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11949 a_578_n57568# a_528_n66# a_314_n57568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11950 GND A6 word438 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11951 a_842_n137656# a_792_n66# a_578_n137656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11952 a_1238_n200# A5 a_974_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11953 a_50_n88240# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11954 a_1898_n39676# a_1848_n66# a_1766_n39676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11955 GND A4 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11956 GND A5 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11957 word589 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11958 a_974_n96760# A6 a_578_n96760# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11959 word122 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11960 word157 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11961 a_1502_n61118# A4 a_1106_n61118# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11962 GND A0 word440 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11963 GND A2 word1002 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11964 word27 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11965 GND A4 word492 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11966 word871 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11967 word652 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11968 word365 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11969 a_1106_n135810# a_1056_n66# a_974_n135810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11970 word736 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11971 a_50_n96192# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11972 a_1898_n115504# a_1848_n66# a_1634_n115504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11973 a_842_n66798# a_792_n66# a_578_n66798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11974 word487 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11975 word218 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11976 word159 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11977 word719 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11978 word1004 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11979 a_182_n56148# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11980 GND A3 word115 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11981 a_1898_n30588# a_1848_n66# a_1766_n30588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11982 GND A0 word338 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11983 a_182_n47770# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11984 a_1502_n38256# A4 a_1238_n38256# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11985 word369 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11986 a_314_n109540# a_264_n66# a_50_n109540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11987 word327 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11988 word386 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11989 a_1502_n60692# A4 a_1106_n60692# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X11990 a_314_n140354# a_264_n66# a_50_n140354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11991 word489 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11992 a_1106_n143762# a_1056_n66# a_842_n143762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11993 a_1634_n135952# a_1584_n66# a_1370_n135952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11994 a_578_n95340# a_528_n66# a_446_n95340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11995 a_314_n131976# a_264_n66# a_50_n131976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11996 GND A6 word645 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11997 GND A3 word662 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X11998 word699 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X11999 word902 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12000 GND A6 word941 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12001 word14 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12002 word329 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12003 word979 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12004 a_974_n132828# A6 a_578_n132828# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12005 word423 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12006 a_1634_n63106# a_1584_n66# a_1370_n63106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12007 a_974_n73188# A6 a_710_n73188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12008 a_314_n117492# a_264_n66# a_50_n117492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12009 a_2294_n14542# A1 a_1898_n14542# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12010 word364 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12011 a_710_n72904# A7 a_446_n72904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12012 a_314_n54160# a_264_n66# a_182_n54160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12013 word110 A0 a_2162_n15820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12014 word945 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12015 a_1238_n84832# A5 a_842_n84832# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12016 a_1634_n104428# a_1584_n66# a_1370_n104428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12017 a_2162_n45924# a_2112_n66# a_2030_n45924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12018 word694 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12019 word425 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12020 a_974_n109966# A6 a_710_n109966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12021 word98 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12022 word635 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12023 word976 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12024 word930 A0 a_2162_n132260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12025 word841 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12026 a_182_n24198# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12027 word166 A0 a_2162_n23772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12028 word915 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12029 word102 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12030 a_578_n63390# a_528_n66# a_314_n63390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12031 a_842_n143478# a_792_n66# a_578_n143478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12032 a_1898_n45498# a_1848_n66# a_1634_n45498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12033 GND A7 word843 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12034 GND A3 word437 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12035 GND A9 word312 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12036 a_2294_n43936# A1 a_1898_n43936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12037 a_1766_n121042# A3 a_1370_n121042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12038 word104 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12039 word303 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12040 word754 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12041 a_710_n40954# A7 a_314_n40954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12042 a_1634_n22778# a_1584_n66# a_1370_n22778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12043 a_1634_n31156# a_1584_n66# a_1370_n31156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12044 word535 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12045 GND A3 word276 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12046 a_1898_n121326# a_1848_n66# a_1766_n121326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12047 word305 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12048 word469 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12049 a_1634_n69638# a_1584_n66# a_1502_n69638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12050 a_710_n87814# A7 a_446_n87814# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12051 word274 A0 a_2162_n39108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12052 a_2030_n69922# A2 a_1634_n69922# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12053 a_314_n69070# a_264_n66# a_182_n69070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12054 GND A7 word779 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12055 a_1106_n127148# a_1056_n66# a_842_n127148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12056 word432 A0 a_2294_n61544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12057 a_2162_n69212# a_2112_n66# a_1898_n69212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12058 GND A6 word824 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12059 GND A5 word94 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12060 a_1238_n21358# A5 a_974_n21358# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12061 word361 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12062 GND A3 word644 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12063 word698 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12064 a_1238_n12980# A5 a_842_n12980# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12065 word370 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12066 a_2030_n107126# A2 a_1766_n107126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12067 word1020 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12068 GND A9 word87 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12069 word207 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12070 a_1634_n60550# a_1584_n66# a_1502_n60550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12071 a_2030_n60834# A2 a_1634_n60834# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12072 a_1238_n68218# A5 a_842_n68218# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12073 GND A5 word582 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12074 word632 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12075 GND A5 word641 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12076 word691 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12077 word210 A0 a_2162_n30020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12078 GND A9 word417 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12079 GND A3 word483 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12080 GND A6 word821 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12081 a_2162_n51746# a_2112_n66# a_2030_n51746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12082 a_2294_n58846# A1 a_1898_n58846# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12083 a_2162_n60124# a_2112_n66# a_1898_n60124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12084 a_2294_n67224# A1 a_2030_n67224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12085 GND A1 word741 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12086 a_1766_n127574# A3 a_1502_n127574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12087 word209 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12088 a_974_n115788# A6 a_710_n115788# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12089 a_1634_n37688# a_1584_n66# a_1502_n37688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12090 a_2030_n37972# A2 a_1634_n37972# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12091 word349 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12092 word882 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12093 a_1898_n136236# a_1848_n66# a_1634_n136236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12094 a_1238_n67792# A5 a_842_n67792# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12095 word575 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12096 word634 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12097 a_2162_n28884# a_2112_n66# a_2030_n28884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12098 word568 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12099 GND A7 word884 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12100 GND A9 word353 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12101 GND A9 word294 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12102 a_2030_n136520# A2 a_1766_n136520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12103 word414 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12104 word795 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12105 GND A5 word199 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12106 word285 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12107 GND A1 word948 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12108 a_1106_n9004# a_1056_n66# a_974_n9004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12109 a_1238_n27890# A5 a_842_n27890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12110 word475 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12111 GND A9 word192 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12112 word615 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12113 a_2030_n144472# A2 a_1634_n144472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12114 a_2294_n26896# A1 a_1898_n26896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12115 a_2162_n129420# a_2112_n66# a_1898_n129420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12116 word183 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12117 word1001 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12118 GND A8 word91 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12119 a_2162_n75034# a_2112_n66# a_1898_n75034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12120 word942 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12121 GND A0 word786 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12122 a_446_n106132# A8 a_50_n106132# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12123 a_1898_n104286# a_1848_n66# a_1634_n104286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12124 a_710_n79152# A7 a_446_n79152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12125 word185 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12126 word671 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12127 a_2162_n137372# a_2112_n66# a_1898_n137372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12128 a_2162_n128994# a_2112_n66# a_2030_n128994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12129 a_1370_n118202# a_1320_n66# a_1106_n118202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12130 a_578_n106416# a_528_n66# a_446_n106416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12131 GND A5 word465 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12132 word721 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12133 a_1238_n74040# A5 a_974_n74040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12134 word673 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12135 word720 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12136 GND A9 word458 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12137 a_2294_n73046# A1 a_2030_n73046# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12138 GND A9 word399 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12139 a_1238_n100452# A5 a_842_n100452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12140 GND A3 word727 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12141 a_710_n39250# A7 a_314_n39250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12142 word250 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12143 word727 a_2376_n66# a_2162_n103434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12144 GND A9 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12145 word267 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12146 a_2030_n43794# A2 a_1766_n43794# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12147 GND A5 word521 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12148 word864 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12149 word981 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12150 a_1898_n142058# a_1848_n66# a_1766_n142058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12151 a_2030_n99032# A2 a_1634_n99032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12152 word729 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12153 a_1238_n138934# A5 a_842_n138934# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12154 a_1898_n133680# a_1848_n66# a_1634_n133680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12155 a_446_n16530# A8 a_182_n16530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12156 a_2162_n43084# a_2112_n66# a_1898_n43084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12157 a_710_n114652# A7 a_314_n114652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12158 word578 A0 a_2162_n82276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12159 GND A8 word137 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12160 GND A8 word196 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12161 word987 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12162 a_578_n135810# a_528_n66# a_314_n135810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12163 a_446_n94204# A8 a_50_n94204# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12164 word514 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12165 a_1898_n119196# a_1848_n66# a_1766_n119196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12166 a_446_n85826# A8 a_50_n85826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12167 a_2294_n132544# A1 a_1898_n132544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12168 a_446_n24482# A8 a_182_n24482# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12169 word507 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12170 GND A1 word16 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12171 GND A7 word823 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12172 GND A3 word993 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12173 GND A1 word989 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12174 a_1106_n6448# a_1056_n66# a_974_n6448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12175 GND A2 word139 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12176 word917 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12177 GND A9 word233 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12178 word993 a_2376_n66# a_2294_n141206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12179 GND A3 word934 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12180 a_2030_n119480# A2 a_1634_n119480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12181 a_2294_n41096# A1 a_2030_n41096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12182 GND A4 word846 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12183 a_578_n143762# a_528_n66# a_314_n143762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12184 a_710_n4602# A7 a_446_n4602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12185 word474 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12186 a_974_n18802# A6 a_578_n18802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12187 GND A3 word832 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12188 a_842_n11702# a_792_n66# a_710_n11702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12189 GND A8 word73 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12190 GND A1 word828 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12191 GND A3 word773 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12192 a_446_n103576# A8 a_50_n103576# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12193 word773 a_2376_n66# a_2294_n109966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12194 a_710_n76596# A7 a_446_n76596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12195 a_1370_n66514# a_1320_n66# a_1238_n66514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12196 word969 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12197 a_2162_n143194# a_2112_n66# a_1898_n143194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12198 word893 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12199 word796 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12200 GND A2 word75 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12201 GND A5 a_1056_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X12202 GND A1 word65 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12203 GND A7 word256 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12204 a_578_n103860# a_528_n66# a_446_n103860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12205 a_1766_n44362# A3 a_1370_n44362# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12206 GND A1 word396 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12207 word21 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12208 GND A9 word499 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12209 a_1502_n124308# A4 a_1106_n124308# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12210 GND A5 word798 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12211 a_1106_n25334# a_1056_n66# a_974_n25334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12212 GND A9 word440 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12213 a_1502_n115930# A4 a_1106_n115930# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12214 a_1106_n16956# a_1056_n66# a_842_n16956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12215 GND A8 word20 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12216 word619 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12217 GND A3 word709 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12218 GND A5 word345 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12219 word249 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12220 word709 a_2376_n66# a_2294_n100878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12221 word1022 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12222 word179 a_2376_n66# a_2162_n25618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12223 word963 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12224 GND A9 word338 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12225 a_1502_n123882# A4 a_1106_n123882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12226 a_710_n120474# A7 a_314_n120474# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12227 a_1370_n34564# a_1320_n66# a_1106_n34564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12228 GND A8 word610 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12229 GND A0 word932 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12230 GND A8 word178 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12231 word667 a_2376_n66# a_2162_n94914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12232 GND A7 word522 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12233 GND A8 word739 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12234 a_50_n143904# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12235 a_1766_n82134# A3 a_1502_n82134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12236 a_2162_n87388# a_2112_n66# a_1898_n87388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12237 word86 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12238 a_1766_n73756# A3 a_1502_n73756# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12239 a_446_n91648# A8 a_50_n91648# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12240 a_1106_n63106# a_1056_n66# a_974_n63106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12241 GND A8 word666 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12242 a_446_n6022# A8 a_182_n6022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12243 a_446_n77164# A8 a_50_n77164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12244 a_1766_n59272# A3 a_1502_n59272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12245 GND A0 word710 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12246 GND A5 word903 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12247 a_974_n24624# A6 a_578_n24624# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12248 a_2294_n85400# A1 a_2030_n85400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12249 word797 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12250 GND A1 word869 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12251 a_1238_n121184# A5 a_842_n121184# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12252 word873 a_2376_n66# a_2294_n124166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12253 a_1370_n72336# a_1320_n66# a_1106_n72336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12254 word571 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12255 GND A0 word262 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12256 word501 a_2376_n66# a_2294_n71342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12257 word875 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12258 a_1370_n121468# a_1320_n66# a_1238_n121468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12259 a_50_n120332# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12260 a_1766_n19370# A3 a_1502_n19370# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12261 GND A7 word297 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12262 a_974_n4176# A6 a_710_n4176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12263 a_50_n111954# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12264 a_1766_n50184# A3 a_1502_n50184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12265 GND A1 word437 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12266 a_1370_n49474# a_1320_n66# a_1238_n49474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12267 GND A5 word780 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12268 GND A7 word627 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12269 word286 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12270 a_578_n23204# a_528_n66# a_446_n23204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12271 word191 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12272 GND A1 word276 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12273 a_1106_n78016# a_1056_n66# a_974_n78016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12274 GND A2 word344 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12275 a_1106_n69638# a_1056_n66# a_842_n69638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12276 GND A4 word992 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12277 word1004 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12278 word620 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12279 GND A4 word933 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12280 a_1370_n40386# a_1320_n66# a_1238_n40386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12281 a_842_n32434# a_792_n66# a_578_n32434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12282 a_974_n39534# A6 a_710_n39534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12283 GND A8 word219 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12284 GND A7 word563 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12285 GND A3 word978 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12286 a_1766_n3324# A3 a_1370_n3324# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12287 a_2162_n8578# a_2112_n66# a_2030_n8578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12288 GND A1 word644 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12289 word902 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12290 word681 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12291 word767 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12292 GND A4 word462 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12293 a_182_n13406# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12294 GND A8 word549 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12295 a_314_n42942# a_264_n66# a_182_n42942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12296 a_1106_n60550# a_1056_n66# a_974_n60550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12297 word883 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12298 word547 a_2376_n66# a_2162_n77874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12299 a_1370_n136378# a_1320_n66# a_1106_n136378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12300 a_446_n3466# A8 a_182_n3466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12301 a_50_n126864# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12302 a_50_n135242# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12303 GND A6 word674 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12304 word391 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12305 a_578_n29736# a_528_n66# a_446_n29736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12306 word703 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12307 word43 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12308 a_50_n91222# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12309 a_842_n70206# a_792_n66# a_578_n70206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12310 word395 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12311 a_974_n77306# A6 a_710_n77306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12312 a_50_n82844# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12313 word325 a_2376_n66# a_2294_n46350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12314 a_1634_n4034# a_1584_n66# a_1370_n4034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12315 a_2294_n5454# A1 a_1898_n5454# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12316 GND A2 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12317 GND A0 word244 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12318 a_1502_n24908# A4 a_1106_n24908# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12319 GND A4 word296 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12320 GND A4 word237 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12321 word955 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12322 a_842_n47344# a_792_n66# a_710_n47344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12323 GND A7 word609 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12324 a_1238_n2614# A5 a_974_n2614# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12325 a_1766_n9856# A3 a_1502_n9856# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12326 a_1898_n11134# a_1848_n66# a_1634_n11134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12327 a_182_n28316# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12328 a_578_n20648# a_528_n66# a_446_n20648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12329 a_50_n103292# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12330 a_842_n100736# a_792_n66# a_578_n100736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12331 a_182_n19938# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12332 a_182_n50752# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12333 a_314_n57852# a_264_n66# a_182_n57852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12334 word131 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12335 a_314_n112522# a_264_n66# a_50_n112522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12336 GND A5 word719 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12337 a_578_n67508# a_528_n66# a_314_n67508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12338 a_1898_n49616# a_1848_n66# a_1634_n49616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12339 word1011 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12340 a_2030_n8152# A2 a_1634_n8152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12341 GND A3 word48 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12342 word58 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12343 a_446_n9998# A8 a_182_n9998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12344 word956 A0 a_2294_n135952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12345 a_974_n36978# A6 a_710_n36978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12346 a_974_n45356# A6 a_710_n45356# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12347 GND A0 word510 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12348 word941 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12349 a_182_n1052# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12350 GND A0 word78 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12351 word749 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12352 a_182_n10850# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12353 a_710_n8294# A7 a_446_n8294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12354 a_50_n97754# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12355 a_842_n85116# a_792_n66# a_710_n85116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12356 a_1370_n84690# a_1320_n66# a_1238_n84690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12357 GND A4 word71 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12358 word229 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12359 a_842_n15394# a_792_n66# a_710_n15394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12360 a_1898_n40528# a_1848_n66# a_1634_n40528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12361 GND A0 word408 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12362 word647 a_2376_n66# a_2162_n92074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12363 word730 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12364 a_182_n57710# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12365 a_50_n132686# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12366 a_50_n141064# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12367 word439 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12368 GND A0 word566 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12369 word734 A0 a_2162_n104428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12370 GND A5 word985 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12371 word561 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12372 word274 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12373 a_314_n141916# a_264_n66# a_50_n141916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12374 word432 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12375 word972 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12376 a_578_n35558# a_528_n66# a_446_n35558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12377 a_1898_n26044# a_1848_n66# a_1766_n26044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12378 GND A6 word283 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12379 a_842_n124024# a_792_n66# a_710_n124024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12380 word278 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12381 word337 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12382 a_182_n65662# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12383 word25 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12384 GND A3 word241 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12385 word493 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12386 a_974_n74750# A6 a_710_n74750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12387 a_314_n127432# a_264_n66# a_50_n127432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12388 a_182_n8010# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12389 a_1634_n1478# a_1584_n66# a_1502_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12390 GND A6 word554 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12391 word1015 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12392 word271 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12393 word716 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12394 a_50_n74182# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12395 a_842_n53166# a_792_n66# a_710_n53166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12396 word332 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12397 a_182_n34138# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12398 GND A4 word608 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12399 a_182_n7584# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12400 a_182_n25760# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12401 a_314_n72052# a_264_n66# a_182_n72052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12402 word236 A0 a_2294_n33712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12403 word214 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12404 a_1370_n99600# a_1320_n66# a_1106_n99600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12405 word393 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12406 a_314_n63674# a_264_n66# a_182_n63674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12407 word231 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12408 word894 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12409 a_1898_n55438# a_1848_n66# a_1766_n55438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12410 word835 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12411 word40 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12412 GND A3 word448 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12413 GND A6 word786 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12414 GND A0 word62 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12415 a_974_n110818# A6 a_710_n110818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12416 word824 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12417 a_974_n42800# A6 a_710_n42800# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12418 word605 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12419 word765 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12420 a_1370_n8152# a_1320_n66# a_1106_n8152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12421 GND A6 word388 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12422 word598 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12423 a_974_n98038# A6 a_578_n98038# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12424 a_2162_n23914# a_2112_n66# a_1898_n23914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12425 a_842_n82560# a_792_n66# a_710_n82560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12426 a_1634_n18234# a_1584_n66# a_1370_n18234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12427 GND A0 word390 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12428 GND A2 word952 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12429 a_1502_n45640# A4 a_1238_n45640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12430 word821 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12431 word661 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12432 word602 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12433 a_50_n89092# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12434 a_842_n68076# a_792_n66# a_578_n68076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12435 a_1898_n93210# a_1848_n66# a_1634_n93210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12436 word168 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12437 word1013 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12438 word431 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12439 a_842_n121468# a_792_n66# a_710_n121468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12440 a_182_n49048# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12441 a_1898_n23488# a_1848_n66# a_1766_n23488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12442 word319 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12443 a_182_n71484# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12444 a_2294_n21926# A1 a_2030_n21926# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12445 a_2294_n30304# A1 a_1898_n30304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12446 a_314_n124876# a_264_n66# a_50_n124876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12447 a_314_n133254# a_264_n66# a_50_n133254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12448 GND A6 word654 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12449 word656 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12450 a_1634_n128852# a_1584_n66# a_1502_n128852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12451 word89 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12452 GND A3 word612 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12453 a_1898_n92784# a_1848_n66# a_1634_n92784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12454 a_1502_n4886# A4 a_1106_n4886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12455 a_1766_n137514# A3 a_1502_n137514# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12456 a_974_n134106# A6 a_578_n134106# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12457 a_1238_n30872# A5 a_842_n30872# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12458 a_1634_n47628# a_1584_n66# a_1502_n47628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12459 a_2030_n47912# A2 a_1766_n47912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12460 word373 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12461 a_1634_n56006# a_1584_n66# a_1502_n56006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12462 word496 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12463 word895 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12464 a_2162_n132402# a_2112_n66# a_2030_n132402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12465 a_314_n47060# a_264_n66# a_182_n47060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12466 a_578_n96192# a_528_n66# a_446_n96192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12467 GND A4 word590 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12468 GND A4 word649 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12469 a_1106_n105138# a_1056_n66# a_842_n105138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12470 GND A4 word64 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12471 a_2162_n47202# a_2112_n66# a_2030_n47202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12472 a_1898_n61260# a_1848_n66# a_1634_n61260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12473 word880 A0 a_2294_n125160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12474 word788 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12475 GND A4 word488 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12476 word543 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12477 a_1502_n82986# A4 a_1238_n82986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12478 a_1502_n91364# A4 a_1238_n91364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12479 a_182_n17098# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12480 GND A0 word44 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12481 word54 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12482 word116 A0 a_2294_n16672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12483 word215 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12484 word865 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12485 word355 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12486 a_578_n56290# a_528_n66# a_314_n56290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12487 a_1898_n38398# a_1848_n66# a_1634_n38398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12488 a_1238_n46208# A5 a_842_n46208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12489 a_1238_n37830# A5 a_974_n37830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12490 GND A3 word387 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12491 GND A9 word262 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12492 a_2294_n45214# A1 a_1898_n45214# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12493 word580 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12494 word113 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12495 a_314_n139786# a_264_n66# a_50_n139786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12496 a_1766_n105564# A3 a_1502_n105564# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12497 word702 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12498 GND A6 word700 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12499 a_710_n42232# A7 a_314_n42232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12500 a_1634_n24056# a_1584_n66# a_1502_n24056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12501 word253 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12502 a_1634_n15678# a_1584_n66# a_1502_n15678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12503 word1012 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12504 GND A5 word266 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12505 a_2162_n100452# a_2112_n66# a_2030_n100452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12506 word727 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12507 a_1238_n45782# A5 a_842_n45782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12508 word478 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12509 word601 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12510 a_2162_n15252# a_2112_n66# a_2030_n15252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12511 word255 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12512 word150 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12513 GND A6 word31 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12514 word382 A0 a_2162_n54444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12515 GND A2 word59 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12516 a_1502_n28600# A4 a_1238_n28600# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12517 word480 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12518 a_1634_n143052# a_1584_n66# a_1502_n143052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12519 a_1106_n142484# a_1056_n66# a_842_n142484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12520 word791 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12521 word318 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12522 a_314_n130698# a_264_n66# a_50_n130698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12523 a_1898_n76170# a_1848_n66# a_1766_n76170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12524 word259 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12525 word690 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12526 a_2294_n104712# A1 a_2030_n104712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12527 word311 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12528 GND A3 word594 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12529 GND A6 word932 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12530 word252 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12531 word379 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12532 a_2294_n74608# A1 a_1898_n74608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12533 a_1766_n143336# A3 a_1370_n143336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12534 GND A1 word793 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12535 word320 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12536 a_1766_n134958# A3 a_1370_n134958# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12537 a_974_n131550# A6 a_578_n131550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12538 a_2294_n13264# A1 a_1898_n13264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12539 a_2030_n53734# A2 a_1634_n53734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12540 a_710_n80004# A7 a_446_n80004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12541 GND A5 word591 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12542 a_2162_n107410# a_2112_n66# a_2030_n107410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12543 GND A5 word532 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12544 word993 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12545 a_710_n10282# A7 a_446_n10282# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12546 a_1238_n83554# A5 a_842_n83554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12547 word685 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12548 GND A6 word771 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12549 a_974_n117066# A6 a_710_n117066# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12550 GND A8 word46 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12551 word376 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12552 a_710_n48764# A7 a_314_n48764# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12553 word648 A0 a_2294_n92216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12554 word832 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12555 a_1898_n129136# a_1848_n66# a_1634_n129136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12556 a_2162_n115362# a_2112_n66# a_2030_n115362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12557 a_2030_n22210# A2 a_1634_n22210# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12558 a_446_n34422# A8 a_182_n34422# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12559 a_1634_n99884# a_1584_n66# a_1370_n99884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12560 GND A7 word834 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12561 GND A7 word893 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12562 a_842_n142200# a_792_n66# a_578_n142200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12563 GND A9 word303 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12564 GND A3 word369 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12565 GND A9 word244 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12566 a_710_n17240# A7 a_446_n17240# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12567 a_2030_n91506# A2 a_1766_n91506# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12568 a_2294_n119622# A1 a_2030_n119622# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12569 a_2030_n30162# A2 a_1766_n30162# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12570 word235 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12571 word95 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12572 a_2030_n21784# A2 a_1634_n21784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12573 a_1238_n29168# A5 a_842_n29168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12574 word416 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12575 GND A8 word143 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12576 a_2162_n82418# a_2112_n66# a_2030_n82418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12577 a_2294_n89518# A1 a_1898_n89518# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12578 word709 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12579 a_1898_n120048# a_1848_n66# a_1634_n120048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12580 a_2162_n21074# a_2112_n66# a_2030_n21074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12581 a_2294_n28174# A1 a_1898_n28174# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12582 a_2030_n68644# A2 a_1766_n68644# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12583 a_710_n86536# A7 a_446_n86536# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12584 word583 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12585 a_2030_n128994# A2 a_1634_n128994# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12586 word843 a_2376_n66# a_2162_n119906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12587 word133 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12588 a_1634_n90796# a_1584_n66# a_1370_n90796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12589 GND A0 word736 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12590 word951 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12591 a_2162_n144756# a_2112_n66# a_2030_n144756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12592 a_1634_n118060# a_1584_n66# a_1370_n118060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12593 word364 A0 a_2294_n51888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12594 word359 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12595 a_2162_n59556# a_2112_n66# a_2030_n59556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12596 a_1634_n140496# a_1584_n66# a_1370_n140496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12597 a_1766_n45924# A3 a_1502_n45924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12598 a_2294_n110534# A1 a_2030_n110534# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12599 GND A5 word85 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12600 word352 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12601 word621 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12602 word694 A0 a_2162_n98748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12603 GND A9 word510 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12604 a_1238_n20080# A5 a_974_n20080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12605 a_2294_n80430# A1 a_1898_n80430# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12606 word630 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12607 GND A9 word78 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12608 GND A5 word415 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12609 word682 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12610 word779 a_2376_n66# a_2162_n110818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12611 word623 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12612 GND A9 word408 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12613 GND A9 word349 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12614 GND A2 word531 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12615 GND A1 word732 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12616 GND A4 word962 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12617 a_1502_n133822# A4 a_1106_n133822# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12618 a_2162_n50468# a_2112_n66# a_2030_n50468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12619 word200 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12620 a_2294_n57568# A1 a_1898_n57568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12621 a_2030_n36694# A2 a_1766_n36694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12622 a_710_n54586# A7 a_314_n54586# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12623 a_1370_n44504# a_1320_n66# a_1106_n44504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12624 GND A5 word471 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12625 word873 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12626 GND A8 word248 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12627 word726 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12628 GND A1 word241 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12629 GND A7 word101 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12630 a_446_n31866# A8 a_182_n31866# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12631 a_1766_n13974# A3 a_1502_n13974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12632 GND A7 word875 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12633 word912 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12634 word528 A0 a_2294_n75176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12635 GND A9 word16 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12636 a_578_n128710# a_528_n66# a_314_n128710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12637 word34 A0 a_2162_n5028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12638 GND A9 word285 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12639 word937 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12640 a_446_n78726# A8 a_50_n78726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12641 a_446_n87104# A8 a_50_n87104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12642 a_1766_n69212# A3 a_1502_n69212# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12643 a_446_n17382# A8 a_182_n17382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12644 word94 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12645 GND A7 word47 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12646 word867 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12647 a_1238_n131124# A5 a_974_n131124# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12648 GND A3 word884 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12649 GND A2 word306 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12650 word808 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12651 GND A9 word183 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12652 word943 a_2376_n66# a_2162_n134106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12653 a_1238_n122746# A5 a_842_n122746# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12654 a_710_n83980# A7 a_446_n83980# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12655 a_2030_n74466# A2 a_1634_n74466# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12656 a_1502_n101872# A4 a_1238_n101872# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12657 a_578_n136662# a_528_n66# a_314_n136662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12658 GND A4 word737 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12659 word848 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12660 a_1370_n12554# a_1320_n66# a_1238_n12554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12661 word992 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12662 a_1370_n131408# a_1320_n66# a_1238_n131408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12663 GND A7 word308 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12664 GND A7 word367 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12665 word933 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12666 GND A1 word837 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12667 a_1766_n60124# A3 a_1502_n60124# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12668 GND A1 word448 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12669 a_2162_n65378# a_2112_n66# a_2030_n65378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12670 GND A9 word65 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12671 a_974_n5738# A6 a_710_n5738# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12672 word978 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12673 a_1106_n32718# a_1056_n66# a_842_n32718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12674 a_1370_n108546# a_1320_n66# a_1106_n108546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12675 a_578_n105138# a_528_n66# a_446_n105138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12676 a_1766_n98606# A3 a_1370_n98606# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12677 word1001 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12678 a_1766_n37262# A3 a_1502_n37262# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12679 word942 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12680 a_1370_n130982# a_1320_n66# a_1238_n130982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12681 word360 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12682 GND A9 word390 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12683 a_1106_n18234# a_1056_n66# a_842_n18234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12684 GND A4 word1003 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12685 word983 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12686 a_2294_n63390# A1 a_1898_n63390# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12687 word129 a_2376_n66# a_2294_n18518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12688 GND A8 word230 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12689 GND A7 word574 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12690 word913 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12691 word972 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12692 a_1238_n137656# A5 a_842_n137656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12693 GND A2 word411 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12694 GND A4 word901 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12695 GND A4 word842 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12696 GND A7 word83 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12697 word287 a_2376_n66# a_2162_n40954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12698 a_1370_n88808# a_1320_n66# a_1106_n88808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12699 a_710_n113374# A7 a_314_n113374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12700 word687 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12701 GND A8 word560 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12702 word953 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12703 word617 a_2376_n66# a_2294_n87814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12704 GND A0 word882 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12705 a_50_n136804# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12706 GND A8 word128 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12707 GND A1 word612 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12708 word919 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12709 a_446_n84548# A8 a_50_n84548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12710 a_1766_n66656# A3 a_1370_n66656# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12711 GND A1 word553 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12712 a_2294_n122888# A1 a_2030_n122888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12713 word776 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12714 GND A1 word121 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12715 GND A6 word57 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12716 GND A6 word312 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12717 GND A8 word616 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12718 a_1106_n5170# a_1056_n66# a_974_n5170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12719 GND A2 word130 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12720 word849 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12721 word925 a_2376_n66# a_2294_n131550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12722 a_710_n3324# A7 a_446_n3324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12723 GND A4 word778 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12724 a_578_n142484# a_528_n66# a_314_n142484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12725 a_842_n10424# a_792_n66# a_710_n10424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12726 GND A2 word618 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12727 GND A3 word823 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12728 a_446_n102298# A8 a_50_n102298# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12729 word823 a_2376_n66# a_2162_n117066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12730 a_842_n48906# a_792_n66# a_710_n48906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12731 word521 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12732 word825 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12733 word728 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12734 word451 a_2376_n66# a_2162_n64242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12735 a_50_n104854# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12736 a_50_n113232# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12737 word243 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12738 GND A1 word328 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12739 GND A5 word789 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12740 a_1502_n123030# A4 a_1106_n123030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12741 GND A5 word730 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12742 a_1106_n24056# a_1056_n66# a_974_n24056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12743 a_2030_n9714# A2 a_1766_n9714# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12744 a_1106_n15678# a_1056_n66# a_842_n15678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12745 a_446_n99458# A8 a_50_n99458# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12746 a_2294_n137798# A1 a_2030_n137798# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12747 a_1502_n484# A4 a_1238_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12748 GND A6 word417 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12749 word954 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12750 word1013 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12751 GND A0 word148 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12752 a_182_n2614# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12753 a_1370_n94630# a_1320_n66# a_1238_n94630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12754 a_710_n9856# A7 a_446_n9856# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12755 GND A4 word141 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12756 a_1898_n910# a_1848_n66# a_1766_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12757 GND A7 word513 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12758 a_842_n16956# a_792_n66# a_710_n16956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12759 a_50_n142626# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12760 word41 a_2376_n66# a_2294_n6022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12761 GND A8 word169 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12762 GND A0 word636 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12763 GND A0 word864 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12764 a_446_n90370# A8 a_50_n90370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12765 word631 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12766 a_1106_n53450# a_1056_n66# a_842_n53450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12767 GND A8 word657 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12768 a_50_n128142# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12769 GND A6 word294 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12770 word348 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12771 a_50_n119764# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12772 GND A5 word835 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12773 word341 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12774 a_974_n23346# A6 a_578_n23346# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12775 GND A2 word659 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12776 word788 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12777 word567 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12778 word786 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12779 a_1370_n71058# a_1320_n66# a_1106_n71058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12780 a_50_n75744# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12781 a_50_n84122# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12782 word343 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12783 word345 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12784 a_1370_n62680# a_1320_n66# a_1106_n62680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12785 word275 a_2376_n66# a_2162_n39250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12786 a_974_n92642# A6 a_578_n92642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12787 GND A0 word194 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12788 word433 a_2376_n66# a_2294_n61686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12789 GND A7 word288 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12790 a_1106_n99884# a_1056_n66# a_974_n99884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12791 a_50_n110676# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12792 word284 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12793 GND A1 word369 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12794 a_1370_n48196# a_1320_n66# a_1238_n48196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12795 a_842_n102014# a_792_n66# a_578_n102014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12796 GND A7 word559 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12797 word758 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12798 a_1766_n87388# A3 a_1502_n87388# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12799 word123 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12800 word182 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12801 a_182_n43652# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12802 GND A3 word86 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12803 a_974_n61118# A6 a_578_n61118# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12804 a_1106_n68360# a_1056_n66# a_842_n68360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12805 GND A6 word399 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12806 word995 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12807 a_578_n91222# a_528_n66# a_446_n91222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12808 a_1106_n90796# a_1056_n66# a_842_n90796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12809 word906 A0 a_2162_n128852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12810 a_974_n38256# A6 a_710_n38256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12811 GND A0 word460 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12812 word23 a_2376_n66# a_2162_n3466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12813 word118 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12814 a_842_n31156# a_792_n66# a_578_n31156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12815 word891 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12816 GND A2 word963 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12817 a_2162_n7300# a_2112_n66# a_2030_n7300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12818 a_974_n60692# A6 a_578_n60692# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12819 word672 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12820 a_182_n12128# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12821 a_50_n99032# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12822 a_578_n59982# a_528_n66# a_314_n59982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12823 GND A4 word453 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12824 a_314_n41664# a_264_n66# a_182_n41664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12825 a_314_n50042# a_264_n66# a_182_n50042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12826 a_842_n69638# a_792_n66# a_578_n69638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12827 word179 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12828 word739 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12829 a_1370_n135100# a_1320_n66# a_1106_n135100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12830 a_446_n2188# A8 a_182_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12831 a_50_n125586# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12832 a_1898_n7868# a_1848_n66# a_1766_n7868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12833 GND A3 word293 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12834 GND A0 word516 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12835 a_314_n134816# a_264_n66# a_50_n134816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12836 GND A6 word665 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12837 word667 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12838 word382 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12839 a_1634_n10708# a_1584_n66# a_1502_n10708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12840 a_974_n20790# A6 a_578_n20790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12841 a_578_n28458# a_528_n66# a_446_n28458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12842 a_842_n108546# a_792_n66# a_578_n108546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12843 a_1238_n40812# A5 a_974_n40812# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12844 a_182_n58562# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12845 a_50_n81566# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12846 GND A3 word132 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12847 a_974_n76028# A6 a_710_n76028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12848 a_2294_n4176# A1 a_1898_n4176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12849 a_578_n97754# a_528_n66# a_446_n97754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12850 GND A2 word24 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12851 a_1502_n23630# A4 a_1106_n23630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12852 a_1502_n32008# A4 a_1106_n32008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12853 GND A2 word738 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12854 GND A4 word228 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12855 a_842_n46066# a_792_n66# a_710_n46066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12856 a_1238_n1336# A5 a_974_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12857 word69 a_2376_n66# a_2294_n9998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12858 GND A7 word600 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12859 word799 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12860 GND A4 word558 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12861 a_182_n18660# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12862 a_182_n27038# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12863 word186 A0 a_2162_n26612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12864 a_1502_n92926# A4 a_1238_n92926# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12865 word1021 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12866 a_314_n56574# a_264_n66# a_182_n56574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12867 a_314_n111244# a_264_n66# a_50_n111244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12868 a_1106_n114652# a_1056_n66# a_974_n114652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12869 word122 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12870 a_578_n66230# a_528_n66# a_314_n66230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12871 GND A6 word440 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12872 a_1634_n106842# a_1584_n66# a_1502_n106842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12873 word501 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12874 word49 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12875 word442 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12876 word1002 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12877 a_842_n137940# a_792_n66# a_578_n137940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12878 a_1502_n78442# A4 a_1106_n78442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12879 word1006 A0 a_2162_n143052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12880 word487 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12881 word124 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12882 a_974_n44078# A6 a_710_n44078# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12883 word555 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12884 word159 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12885 word932 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12886 GND A5 word336 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12887 word740 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12888 a_1238_n55722# A5 a_974_n55722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12889 GND A4 word494 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12890 word548 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12891 a_50_n96476# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12892 word220 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12893 a_1634_n94914# a_1584_n66# a_1370_n94914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12894 GND A0 word340 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12895 a_1502_n38540# A4 a_1238_n38540# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12896 word552 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12897 word771 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12898 GND A4 word333 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12899 a_1502_n60976# A4 a_1106_n60976# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12900 a_314_n140638# a_264_n66# a_50_n140638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12901 a_1634_n144614# a_1584_n66# a_1370_n144614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12902 word26 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12903 a_1898_n86110# a_1848_n66# a_1634_n86110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12904 word710 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12905 word423 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12906 word364 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12907 word381 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12908 a_578_n34280# a_528_n66# a_446_n34280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12909 GND A6 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12910 a_842_n105990# a_792_n66# a_578_n105990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12911 a_182_n64384# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12912 a_1502_n46492# A4 a_1238_n46492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12913 a_314_n126154# a_264_n66# a_50_n126154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12914 a_2030_n132402# A2 a_1766_n132402# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12915 a_314_n117776# a_264_n66# a_50_n117776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12916 GND A6 word545 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12917 a_1898_n94062# a_1848_n66# a_1766_n94062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12918 a_710_n11844# A7 a_446_n11844# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12919 a_1502_n6164# A4 a_1106_n6164# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12920 word707 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12921 VDD A5 a_1056_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X12922 a_1634_n62964# a_1584_n66# a_1370_n62964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12923 word843 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12924 a_2162_n116924# a_2112_n66# a_1898_n116924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12925 a_314_n62396# a_264_n66# a_182_n62396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12926 word163 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12927 a_1898_n54160# a_1848_n66# a_1634_n54160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12928 a_1634_n112664# a_1584_n66# a_1370_n112664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12929 word535 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12930 word830 A0 a_2162_n118060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12931 GND A3 word439 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12932 word988 A0 a_2294_n140496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12933 GND A6 word777 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12934 word63 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12935 word97 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12936 word224 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12937 a_1766_n121326# A3 a_1370_n121326# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12938 word651 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12939 word469 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12940 a_1634_n31440# a_1584_n66# a_1370_n31440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12941 a_2030_n40102# A2 a_1634_n40102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12942 word305 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12943 word486 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12944 a_2030_n100452# A2 a_1766_n100452# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12945 a_1238_n39108# A5 a_974_n39108# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12946 GND A3 word337 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12947 a_1898_n121610# a_1848_n66# a_1766_n121610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12948 GND A3 word278 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12949 a_2030_n138934# A2 a_1766_n138934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12950 a_2162_n22636# a_2112_n66# a_1898_n22636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12951 word203 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12952 a_2294_n29736# A1 a_2030_n29736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12953 word221 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12954 word361 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12955 word434 A0 a_2162_n61828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12956 word962 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12957 a_1238_n38682# A5 a_974_n38682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12958 word370 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12959 a_2162_n91932# a_2112_n66# a_1898_n91932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12960 GND A5 word155 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12961 word422 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12962 a_1634_n86252# a_1584_n66# a_1370_n86252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12963 word691 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12964 a_446_n12412# A8 a_182_n12412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12965 a_1238_n30020# A5 a_842_n30020# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12966 word363 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12967 a_842_n120190# a_792_n66# a_710_n120190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12968 GND A7 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12969 word332 A0 a_2294_n47344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12970 a_2030_n107410# A2 a_1766_n107410# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12971 GND A9 word148 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12972 GND A3 word214 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12973 word741 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12974 GND A9 word89 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12975 a_1106_n135384# a_1056_n66# a_974_n135384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12976 a_2294_n20648# A1 a_2030_n20648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12977 a_1898_n69070# a_1848_n66# a_1766_n69070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12978 a_314_n123598# a_264_n66# a_50_n123598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12979 GND A5 word643 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12980 word647 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12981 word693 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12982 word426 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12983 GND A5 word211 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12984 GND A3 word544 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12985 GND A5 word152 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12986 a_1766_n127858# A3 a_1502_n127858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12987 a_2030_n55012# A2 a_1766_n55012# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12988 a_2030_n115362# A2 a_1634_n115362# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12989 GND A5 word541 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12990 a_2030_n106984# A2 a_1766_n106984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12991 word1019 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12992 GND A4 word640 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12993 word884 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12994 a_2162_n131124# a_2112_n66# a_2030_n131124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X12995 a_2162_n122746# a_2112_n66# a_1898_n122746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12996 a_1238_n76454# A5 a_974_n76454# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12997 a_2162_n37546# a_2112_n66# a_1898_n37546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X12998 word737 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X12999 a_1766_n23914# A3 a_1502_n23914# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13000 word326 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13001 word598 A0 a_2162_n85116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13002 word407 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13003 GND A9 word355 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13004 word45 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13005 word475 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13006 word534 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13007 a_2030_n15110# A2 a_1634_n15110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13008 GND A5 word260 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13009 a_446_n27322# A8 a_182_n27322# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13010 a_446_n18944# A8 a_182_n18944# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13011 GND A1 word36 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13012 GND A9 word253 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13013 GND A9 word194 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13014 a_2030_n84406# A2 a_1766_n84406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13015 a_2030_n144756# A2 a_1634_n144756# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13016 a_2294_n35558# A1 a_2030_n35558# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13017 a_2030_n23062# A2 a_1766_n23062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13018 word185 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13019 GND A5 word257 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13020 GND A8 word93 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13021 word1003 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13022 word718 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13023 a_2162_n66940# a_2112_n66# a_1898_n66940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13024 a_446_n106416# A8 a_50_n106416# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13025 a_1898_n104570# a_1848_n66# a_1634_n104570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13026 a_1238_n109824# A5 a_974_n109824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13027 a_710_n79436# A7 a_446_n79436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13028 word592 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13029 a_1106_n8862# a_1056_n66# a_974_n8862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13030 word673 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13031 a_710_n18092# A7 a_446_n18092# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13032 GND A6 word22 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13033 word491 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13034 a_1634_n83696# a_1584_n66# a_1502_n83696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13035 GND A2 word50 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13036 word901 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13037 GND A8 word581 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13038 word314 A0 a_2162_n44788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13039 word723 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13040 a_1370_n140922# a_1320_n66# a_1238_n140922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13041 a_1634_n133396# a_1584_n66# a_1502_n133396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13042 word250 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13043 a_1766_n38824# A3 a_1370_n38824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13044 word41 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13045 a_2162_n74892# a_2112_n66# a_1898_n74892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13046 word302 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13047 GND A6 word923 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13048 GND A9 word460 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13049 GND A7 word776 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13050 a_1766_n142058# A3 a_1502_n142058# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13051 GND A1 word784 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13052 a_1238_n100736# A5 a_842_n100736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13053 word729 a_2376_n66# a_2294_n103718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13054 a_2030_n52456# A2 a_1766_n52456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13055 GND A5 word523 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13056 word427 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13057 a_1238_n73898# A5 a_974_n73898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13058 GND A2 word481 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13059 a_1238_n82276# A5 a_842_n82276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13060 a_2030_n99316# A2 a_1634_n99316# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13061 a_1766_n119196# A3 a_1502_n119196# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13062 a_710_n123314# A7 a_314_n123314# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13063 GND A1 word293 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13064 a_710_n114936# A7 a_314_n114936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13065 a_710_n47486# A7 a_314_n47486# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13066 GND A8 word37 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13067 word507 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13068 GND A8 word198 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13069 word580 A0 a_2294_n82560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13070 word764 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13071 a_2162_n114084# a_2112_n66# a_2030_n114084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13072 word266 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13073 GND A8 word139 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13074 word989 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13075 a_2294_n141206# A1 a_2030_n141206# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13076 word846 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13077 a_446_n33144# A8 a_182_n33144# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13078 a_446_n24766# A8 a_182_n24766# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13079 GND A1 word132 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13080 word509 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13081 GND A7 word825 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13082 GND A8 word686 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13083 word478 A0 a_2162_n68076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13084 GND A9 word235 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13085 word887 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13086 a_2030_n90228# A2 a_1634_n90228# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13087 GND A8 word756 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13088 a_2294_n118344# A1 a_2030_n118344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13089 GND A3 word690 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13090 a_2294_n109966# A1 a_1898_n109966# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13091 GND A7 word56 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13092 a_2294_n88240# A1 a_1898_n88240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13093 GND A8 word75 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13094 a_2162_n81140# a_2112_n66# a_2030_n81140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13095 word817 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13096 GND A9 word133 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13097 word893 a_2376_n66# a_2294_n127006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13098 GND A1 word889 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13099 GND A3 word834 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13100 GND A2 word256 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13101 a_710_n85258# A7 a_446_n85258# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13102 a_446_n103860# A8 a_50_n103860# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13103 word633 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13104 a_578_n129562# a_528_n66# a_314_n129562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13105 GND A4 word746 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13106 a_710_n76880# A7 a_446_n76880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13107 a_2030_n67366# A2 a_1634_n67366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13108 word591 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13109 word798 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13110 GND A7 word317 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13111 GND A7 word258 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13112 a_974_n7016# A6 a_710_n7016# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13113 a_2162_n49900# a_2112_n66# a_1898_n49900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13114 a_1766_n53024# A3 a_1370_n53024# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13115 a_2294_n96192# A1 a_1898_n96192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13116 word23 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13117 a_2294_n100878# A1 a_1898_n100878# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13118 a_1106_n25618# a_1056_n66# a_974_n25618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13119 word892 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13120 word614 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13121 GND A2 word522 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13122 GND A9 word340 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13123 GND A5 word856 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13124 a_2030_n96760# A2 a_1634_n96760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13125 a_1502_n132544# A4 a_1106_n132544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13126 a_710_n120758# A7 a_314_n120758# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13127 GND A8 word19 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13128 a_1370_n34848# a_1320_n66# a_1106_n34848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13129 word366 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13130 GND A8 word239 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13131 a_2162_n96050# a_2112_n66# a_2030_n96050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13132 GND A7 word524 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13133 GND A0 word934 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13134 GND A8 word180 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13135 a_1766_n82418# A3 a_1502_n82418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13136 word237 a_2376_n66# a_2294_n33854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13137 GND A7 word92 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13138 a_1502_n109682# A4 a_1238_n109682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13139 a_1766_n21074# A3 a_1370_n21074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13140 GND A1 word232 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13141 word696 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13142 a_446_n30588# A8 a_182_n30588# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13143 GND A1 word173 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13144 GND A9 word7 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13145 a_1370_n139218# a_1320_n66# a_1238_n139218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13146 a_1502_n101020# A4 a_1238_n101020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13147 GND A0 word832 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13148 a_446_n6306# A8 a_182_n6306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13149 a_50_n129704# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13150 word869 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13151 a_446_n77448# A8 a_50_n77448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13152 a_1766_n59556# A3 a_1502_n59556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13153 GND A8 word738 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13154 a_2294_n124166# A1 a_2030_n124166# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13155 a_1766_n81992# A3 a_1502_n81992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13156 GND A5 word905 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13157 word69 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13158 a_2162_n2330# a_2112_n66# a_1898_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13159 a_974_n24908# A6 a_578_n24908# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13160 GND A7 word38 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13161 GND A6 word262 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13162 a_1106_n71342# a_1056_n66# a_842_n71342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13163 word799 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13164 word858 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13165 a_1238_n121468# A5 a_842_n121468# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13166 GND A2 word297 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13167 a_1106_n62964# a_1056_n66# a_974_n62964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13168 a_2030_n73188# A2 a_1766_n73188# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13169 a_1370_n138792# a_1320_n66# a_1238_n138792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13170 word875 a_2376_n66# a_2162_n124450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13171 a_578_n135384# a_528_n66# a_314_n135384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13172 word415 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13173 a_1370_n72620# a_1320_n66# a_1106_n72620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13174 a_1502_n100594# A4 a_1238_n100594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13175 GND A5 word669 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13176 word56 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13177 word573 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13178 word503 a_2376_n66# a_2162_n71626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13179 GND A7 word358 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13180 GND A2 word627 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13181 GND A5 word961 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13182 a_1370_n130130# a_1320_n66# a_1238_n130130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13183 a_50_n120616# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13184 a_2162_n64100# a_2112_n66# a_2030_n64100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13185 GND A7 word299 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13186 GND A1 word769 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13187 a_974_n4460# A6 a_710_n4460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13188 word71 a_2376_n66# a_2162_n10282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13189 a_1766_n50468# A3 a_1502_n50468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13190 a_1370_n49758# a_1320_n66# a_1238_n49758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13191 a_1370_n58136# a_1320_n66# a_1238_n58136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13192 a_1370_n80572# a_1320_n66# a_1106_n80572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13193 GND A7 word629 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13194 word401 a_2376_n66# a_2294_n57142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13195 a_1370_n107268# a_1320_n66# a_1106_n107268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13196 a_50_n106132# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13197 a_1766_n88950# A3 a_1370_n88950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13198 GND A1 word337 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13199 GND A2 word563 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13200 GND A4 word994 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13201 GND A2 word504 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13202 GND A4 word935 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13203 a_842_n32718# a_792_n66# a_578_n32718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13204 a_974_n39818# A6 a_710_n39818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13205 word190 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13206 a_1370_n40670# a_1320_n66# a_1238_n40670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13207 GND A7 word565 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13208 GND A3 word980 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13209 word904 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13210 a_1238_n128000# A5 a_974_n128000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13211 GND A0 word98 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13212 a_578_n69922# a_528_n66# a_314_n69922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13213 GND A2 word402 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13214 a_1106_n77874# a_1056_n66# a_974_n77874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13215 a_2030_n88098# A2 a_1634_n88098# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13216 a_710_n112096# A7 a_314_n112096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13217 GND A4 word833 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13218 word944 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13219 a_314_n51604# a_264_n66# a_182_n51604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13220 a_1370_n26186# a_1320_n66# a_1106_n26186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13221 a_1370_n145040# a_1320_n66# a_1106_n145040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13222 word885 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13223 a_842_n18234# a_792_n66# a_710_n18234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13224 GND A8 word119 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13225 GND A0 word814 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13226 a_50_n135526# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13227 GND A1 word544 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13228 GND A0 word586 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13229 a_446_n3750# A8 a_182_n3750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13230 a_446_n83270# A8 a_50_n83270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13231 a_1766_n57000# A3 a_1370_n57000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13232 word766 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13233 a_182_n21642# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13234 a_1370_n95482# a_1320_n66# a_1238_n95482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13235 GND A6 word303 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13236 GND A8 word607 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13237 a_842_n140922# a_792_n66# a_578_n140922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13238 word806 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13239 a_710_n2046# A7 a_446_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13240 a_182_n68502# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13241 a_50_n91506# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13242 a_578_n60834# a_528_n66# a_314_n60834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13243 a_1898_n42942# a_1848_n66# a_1634_n42942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13244 a_1634_n4318# a_1584_n66# a_1370_n4318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13245 GND A2 word609 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13246 GND A2 word867 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13247 GND A2 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13248 a_1898_n89802# a_1848_n66# a_1766_n89802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13249 word736 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13250 GND A2 word808 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13251 word517 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13252 a_50_n77022# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13253 GND A4 word298 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13254 a_842_n47628# a_792_n66# a_710_n47628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13255 a_1370_n113090# a_1320_n66# a_1238_n113090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13256 a_1898_n11418# a_1848_n66# a_1634_n11418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13257 word383 a_2376_n66# a_2162_n54586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13258 a_314_n66514# a_264_n66# a_182_n66514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13259 a_50_n103576# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13260 a_1634_n3892# a_1584_n66# a_1370_n3892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13261 GND A4 word196 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13262 GND A4 word137 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13263 a_1502_n41522# A4 a_1106_n41522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13264 a_314_n112806# a_264_n66# a_50_n112806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13265 GND A0 word978 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13266 word767 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13267 a_1106_n14400# a_1056_n66# a_842_n14400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13268 word60 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13269 a_446_n98180# A8 a_50_n98180# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13270 a_1898_n80714# a_1848_n66# a_1766_n80714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13271 GND A0 word632 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13272 a_2030_n8436# A2 a_1634_n8436# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13273 a_1898_n10992# a_1848_n66# a_1634_n10992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13274 a_182_n36552# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13275 word229 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13276 GND A6 word408 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13277 word945 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13278 word810 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13279 GND A0 word80 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13280 a_1898_n57852# a_1848_n66# a_1766_n57852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13281 GND A6 word566 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13282 word911 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13283 a_182_n1336# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13284 a_710_n8578# A7 a_446_n8578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13285 word561 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13286 word985 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13287 GND A4 word73 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13288 word127 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13289 GND A0 word410 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13290 word649 a_2376_n66# a_2294_n92358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13291 a_842_n15678# a_792_n66# a_710_n15678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13292 a_50_n141348# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13293 GND A0 word568 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13294 GND A1 word585 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13295 word703 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13296 word622 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13297 word841 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13298 GND A2 word913 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13299 a_50_n132970# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13300 a_1766_n71200# A3 a_1370_n71200# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13301 word493 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13302 word434 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13303 word866 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13304 word807 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13305 word129 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13306 word974 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13307 GND A6 word285 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13308 a_842_n84974# a_792_n66# a_710_n84974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13309 a_842_n124308# a_792_n66# a_710_n124308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13310 a_50_n118486# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13311 a_1898_n9146# a_1848_n66# a_1634_n9146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13312 a_1898_n17950# a_1848_n66# a_1634_n17950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13313 word339 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13314 GND A0 word466 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13315 word847 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13316 GND A3 word243 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13317 word280 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13318 a_1502_n56432# A4 a_1238_n56432# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13319 word497 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13320 word792 A0 a_2294_n112664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13321 a_182_n65946# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13322 a_314_n127716# a_264_n66# a_50_n127716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13323 word332 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13324 a_974_n22068# A6 a_578_n22068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13325 GND A2 word650 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13326 word273 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13327 GND A6 word183 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13328 word777 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13329 GND A2 word849 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13330 a_842_n123882# a_792_n66# a_710_n123882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13331 a_50_n74466# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13332 a_842_n53450# a_792_n66# a_710_n53450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13333 word334 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13334 a_578_n99032# a_528_n66# a_446_n99032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13335 a_974_n91364# A6 a_578_n91364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13336 GND A6 word671 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13337 GND A4 word610 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13338 GND A2 word747 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13339 a_182_n7868# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13340 a_314_n72336# a_264_n66# a_182_n72336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13341 a_314_n63958# a_264_n66# a_182_n63958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13342 a_1634_n122604# a_1584_n66# a_1370_n122604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13343 word174 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13344 word605 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13345 word695 a_2376_n66# a_2162_n98890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13346 GND A7 word550 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13347 word749 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13348 a_2030_n5880# A2 a_1634_n5880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13349 word167 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13350 word136 A0 a_2294_n19512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13351 word114 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13352 a_182_n33996# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13353 a_182_n42374# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13354 a_314_n49474# a_264_n66# a_182_n49474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13355 a_1502_n24482# A4 a_1106_n24482# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13356 a_1106_n107552# a_1056_n66# a_842_n107552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13357 a_1370_n8436# a_1320_n66# a_1106_n8436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13358 a_578_n59130# a_528_n66# a_314_n59130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13359 GND A6 word390 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13360 word392 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13361 word451 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13362 a_842_n139218# a_792_n66# a_578_n139218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13363 a_1898_n63674# a_1848_n66# a_1634_n63674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13364 word661 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13365 word602 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13366 word109 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13367 a_2030_n18802# A2 a_1766_n18802# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13368 word431 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13369 word882 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13370 word663 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13371 GND A2 word954 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13372 a_578_n67082# a_528_n66# a_314_n67082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13373 a_1634_n40954# a_1584_n66# a_1370_n40954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13374 word604 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13375 a_842_n138792# a_792_n66# a_578_n138792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13376 a_50_n89376# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13377 word72 A0 a_2294_n10424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13378 a_1238_n48622# A5 a_842_n48622# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13379 GND A4 word385 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13380 a_314_n40386# a_264_n66# a_182_n40386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13381 a_842_n68360# a_792_n66# a_578_n68360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13382 word170 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13383 word1015 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13384 a_842_n90796# a_792_n66# a_710_n90796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13385 word597 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13386 a_1634_n87814# a_1584_n66# a_1502_n87814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13387 a_974_n97896# A6 a_578_n97896# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13388 a_1898_n6590# a_1848_n66# a_1634_n6590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13389 word380 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13390 a_1106_n145324# a_1056_n66# a_842_n145324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13391 a_182_n71768# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13392 word279 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13393 a_314_n133538# a_264_n66# a_50_n133538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13394 word658 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13395 word373 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13396 word314 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13397 a_578_n27180# a_528_n66# a_446_n27180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13398 GND A5 word281 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13399 word226 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13400 a_842_n107268# a_792_n66# a_578_n107268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13401 GND A5 word222 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13402 a_182_n57284# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13403 GND A3 word182 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13404 a_2030_n125302# A2 a_1766_n125302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13405 a_50_n80288# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13406 a_2294_n16104# A1 a_2030_n16104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13407 word375 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13408 a_314_n119054# a_264_n66# a_50_n119054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13409 word498 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13410 a_710_n13122# A7 a_446_n13122# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13411 a_578_n96476# a_528_n66# a_446_n96476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13412 GND A3 word611 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13413 word215 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13414 a_974_n133964# A6 a_578_n133964# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13415 a_1766_n7300# A3 a_1370_n7300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13416 word477 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13417 a_2162_n118202# a_2112_n66# a_1898_n118202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13418 word790 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13419 a_1634_n55864# a_1584_n66# a_1502_n55864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13420 GND A4 word549 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13421 a_1502_n91648# A4 a_1238_n91648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13422 word118 A0 a_2162_n16956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13423 GND A4 word490 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13424 a_314_n55296# a_264_n66# a_182_n55296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13425 a_842_n145040# a_792_n66# a_578_n145040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13426 a_1106_n104996# a_1056_n66# a_842_n104996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13427 word702 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13428 word433 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13429 word492 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13430 word106 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13431 GND A3 word389 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13432 word938 A0 a_2162_n133396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13433 word115 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13434 a_1502_n68786# A4 a_1106_n68786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13435 word478 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13436 word419 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13437 a_1766_n114226# A3 a_1502_n114226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13438 word255 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13439 a_710_n42516# A7 a_314_n42516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13440 word150 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13441 a_1634_n24340# a_1584_n66# a_1502_n24340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13442 GND A5 word327 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13443 GND A5 word386 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13444 word923 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13445 word864 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13446 GND A2 word995 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13447 word645 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13448 word729 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13449 a_50_n95198# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13450 a_1898_n114510# a_1848_n66# a_1766_n114510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13451 word603 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13452 word638 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13453 word311 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13454 a_974_n110392# A6 a_710_n110392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13455 word912 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13456 word384 A0 a_2294_n54728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13457 word379 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13458 a_1106_n142768# a_1056_n66# a_842_n142768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13459 word793 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13460 word895 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13461 a_1898_n122462# a_1848_n66# a_1634_n122462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13462 word372 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13463 a_1634_n79152# a_1584_n66# a_1502_n79152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13464 word313 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13465 GND A6 word934 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13466 a_1766_n143620# A3 a_1370_n143620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13467 GND A3 word164 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13468 GND A7 word787 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13469 GND A7 word846 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13470 GND A9 word98 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13471 a_2030_n131124# A2 a_1634_n131124# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13472 a_314_n116498# a_264_n66# a_50_n116498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13473 GND A5 word593 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13474 a_710_n10566# A7 a_446_n10566# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13475 a_1238_n83838# A5 a_842_n83838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13476 a_1238_n92216# A5 a_974_n92216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13477 GND A6 word773 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13478 a_1238_n22494# A5 a_974_n22494# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13479 a_2162_n44930# a_2112_n66# a_2030_n44930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13480 a_2162_n53308# a_2112_n66# a_1898_n53308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13481 a_2294_n91222# A1 a_2030_n91222# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13482 a_974_n117350# A6 a_710_n117350# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13483 word378 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13484 a_2030_n108262# A2 a_1634_n108262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13485 a_1634_n70064# a_1584_n66# a_1502_n70064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13486 word577 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13487 word893 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13488 word969 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13489 word746 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13490 word834 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13491 a_1898_n129420# a_1848_n66# a_1634_n129420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13492 word218 A0 a_2162_n31156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13493 word154 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13494 a_1634_n111386# a_1584_n66# a_1502_n111386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13495 a_446_n34706# A8 a_182_n34706# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13496 word95 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13497 a_1766_n16814# A3 a_1370_n16814# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13498 a_2162_n52882# a_2112_n66# a_2030_n52882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13499 a_2294_n59982# A1 a_1898_n59982# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13500 word548 A0 a_2294_n78016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13501 GND A9 word305 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13502 GND A9 word36 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13503 a_2294_n51320# A1 a_2030_n51320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13504 a_1766_n111670# A3 a_1370_n111670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13505 word583 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13506 word642 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13507 a_1898_n137372# a_1848_n66# a_1766_n137372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13508 word418 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13509 GND A7 word67 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13510 GND A9 word203 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13511 GND A7 word892 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13512 a_578_n139502# a_528_n66# a_314_n139502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13513 a_710_n86820# A7 a_446_n86820# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13514 a_1502_n104712# A4 a_1106_n104712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13515 GND A9 word361 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13516 a_2030_n137656# A2 a_1634_n137656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13517 a_2162_n12980# a_2112_n66# a_2030_n12980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13518 word135 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13519 a_2294_n50894# A1 a_1898_n50894# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13520 word953 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13521 GND A5 word207 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13522 a_2162_n68218# a_2112_n66# a_1898_n68218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13523 word111 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13524 a_1634_n140780# a_1584_n66# a_1370_n140780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13525 word483 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13526 GND A1 word956 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13527 a_446_n11134# A8 a_182_n11134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13528 word354 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13529 a_1634_n76596# a_1584_n66# a_1370_n76596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13530 word623 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13531 GND A8 word531 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13532 word264 A0 a_2294_n37688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13533 GND A9 word80 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13534 word684 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13535 a_1634_n126296# a_1584_n66# a_1370_n126296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13536 a_578_n130414# a_528_n66# a_314_n130414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13537 word625 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13538 GND A3 word535 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13539 GND A9 word410 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13540 a_2294_n66230# A1 a_2030_n66230# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13541 a_1238_n102014# A5 a_842_n102014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13542 GND A6 word814 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13543 a_578_n107552# a_528_n66# a_446_n107552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13544 a_2030_n114084# A2 a_1766_n114084# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13545 a_2030_n36978# A2 a_1766_n36978# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13546 GND A5 word473 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13547 word377 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13548 GND A5 word414 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13549 a_1238_n75176# A5 a_974_n75176# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13550 word875 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13551 a_2162_n121468# a_2112_n66# a_1898_n121468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13552 a_1238_n66798# A5 a_842_n66798# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13553 word728 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13554 GND A9 word466 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13555 a_2162_n36268# a_2112_n66# a_1898_n36268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13556 GND A7 word103 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13557 a_710_n116214# A7 a_314_n116214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13558 GND A9 word407 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13559 a_1502_n119622# A4 a_1238_n119622# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13560 a_2162_n27890# a_2112_n66# a_2030_n27890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13561 a_2294_n74182# A1 a_2030_n74182# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13562 word457 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13563 word530 A0 a_2162_n75460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13564 GND A9 word18 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13565 GND A0 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13566 word939 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13567 word796 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13568 a_710_n342# A7 a_446_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13569 a_1766_n91932# A3 a_1502_n91932# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13570 a_1898_n143194# a_1848_n66# a_1634_n143194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13571 a_2294_n125728# A1 a_1898_n125728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13572 a_446_n17666# A8 a_182_n17666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13573 a_446_n26044# A8 a_182_n26044# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13574 word155 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13575 a_1106_n8010# a_1056_n66# a_974_n8010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13576 a_1238_n131408# A5 a_974_n131408# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13577 GND A9 word185 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13578 word837 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13579 a_578_n145324# a_528_n66# a_314_n145324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13580 a_2294_n34280# A1 a_2030_n34280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13581 a_2030_n83128# A2 a_1634_n83128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13582 a_2030_n143478# A2 a_1766_n143478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13583 a_578_n136946# a_528_n66# a_314_n136946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13584 a_1502_n110534# A4 a_1238_n110534# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13585 a_1370_n21216# a_1320_n66# a_1238_n21216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13586 a_446_n86962# A8 a_50_n86962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13587 word994 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13588 a_1370_n12838# a_1320_n66# a_1238_n12838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13589 GND A8 word84 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13590 word935 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13591 word141 a_2376_n66# a_2294_n20222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13592 word152 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13593 a_446_n105138# A8 a_50_n105138# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13594 a_1106_n7584# a_1056_n66# a_974_n7584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13595 a_710_n78158# A7 a_446_n78158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13596 word1001 a_2376_n66# a_2294_n142342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13597 GND A1 word997 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13598 a_1238_n130982# A5 a_974_n130982# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13599 GND A1 word77 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13600 GND A6 word13 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13601 word541 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13602 a_1370_n90512# a_1320_n66# a_1106_n90512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13603 word980 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13604 GND A8 word572 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13605 a_2162_n136378# a_2112_n66# a_1898_n136378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13606 a_1370_n117208# a_1320_n66# a_1106_n117208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13607 GND A7 word267 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13608 a_1370_n108830# a_1320_n66# a_1106_n108830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13609 word1003 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13610 GND A1 word348 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13611 a_1766_n37546# A3 a_1502_n37546# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13612 GND A4 word1005 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13613 GND A3 word720 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13614 GND A2 word83 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13615 word842 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13616 a_1370_n116782# a_1320_n66# a_1106_n116782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13617 a_578_n104996# a_528_n66# a_446_n104996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13618 GND A5 word514 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13619 word974 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13620 GND A2 word472 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13621 a_1106_n87814# a_1056_n66# a_842_n87814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13622 a_2030_n98038# A2 a_1766_n98038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13623 GND A9 word507 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13624 a_1238_n137940# A5 a_842_n137940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13625 GND A4 word903 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13626 a_2162_n42090# a_2112_n66# a_1898_n42090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13627 a_2294_n49190# A1 a_2030_n49190# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13628 a_710_n113658# A7 a_314_n113658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13629 a_710_n122036# A7 a_314_n122036# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13630 GND A1 word284 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13631 GND A8 word28 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13632 word955 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13633 a_1370_n36126# a_1320_n66# a_1106_n36126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13634 GND A0 word884 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13635 word316 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13636 GND A8 word130 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13637 GND A8 word189 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13638 a_446_n93210# A8 a_50_n93210# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13639 a_1766_n75318# A3 a_1370_n75318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13640 word187 a_2376_n66# a_2162_n26754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13641 a_1766_n66940# A3 a_1370_n66940# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13642 a_2294_n131550# A1 a_1898_n131550# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13643 word778 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13644 a_446_n23488# A8 a_182_n23488# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13645 word500 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13646 GND A1 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13647 GND A6 word59 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13648 GND A8 word677 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13649 word1011 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13650 GND A8 word618 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13651 GND A8 word747 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13652 word819 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13653 GND A4 word780 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13654 a_578_n142768# a_528_n66# a_314_n142768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13655 a_710_n3608# A7 a_446_n3608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13656 a_2294_n108688# A1 a_1898_n108688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13657 a_446_n92784# A8 a_50_n92784# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13658 a_842_n10708# a_792_n66# a_710_n10708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13659 GND A1 word880 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13660 a_2030_n66088# A2 a_1766_n66088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13661 word825 a_2376_n66# a_2294_n117350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13662 a_578_n128284# a_528_n66# a_314_n128284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13663 word789 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13664 word523 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13665 GND A0 word718 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13666 GND A5 word911 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13667 word730 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13668 word453 a_2376_n66# a_2294_n64526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13669 a_50_n113516# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13670 GND A1 word389 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13671 a_1766_n34990# A3 a_1370_n34990# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13672 a_1766_n43368# A3 a_1370_n43368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13673 a_1106_n24340# a_1056_n66# a_974_n24340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13674 GND A6 word148 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13675 a_1502_n768# A4 a_1238_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13676 word1015 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13677 GND A2 word513 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13678 GND A2 word712 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13679 GND A5 word847 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13680 word631 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13681 a_1502_n122888# A4 a_1106_n122888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13682 a_1106_n32292# a_1056_n66# a_842_n32292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13683 GND A4 word143 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13684 word43 a_2376_n66# a_2162_n6306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13685 a_1106_n79152# a_1056_n66# a_974_n79152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13686 GND A7 word515 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13687 a_1238_n129278# A5 a_974_n129278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13688 a_50_n142910# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13689 a_974_n63532# A6 a_578_n63532# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13690 word936 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13691 word877 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13692 a_314_n44504# a_264_n66# a_182_n44504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13693 GND A1 word164 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13694 word894 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13695 GND A4 word46 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13696 GND A0 word536 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13697 GND A0 word764 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13698 GND A8 word659 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13699 a_446_n5028# A8 a_182_n5028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13700 a_50_n128426# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13701 a_446_n76170# A8 a_50_n76170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13702 GND A7 word571 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13703 GND A6 a_792_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X13704 word567 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13705 GND A1 word652 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13706 word862 A0 a_2162_n122604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13707 word343 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13708 a_182_n14542# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13709 a_974_n23630# A6 a_578_n23630# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13710 GND A8 word557 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13711 a_578_n62112# a_528_n66# a_314_n62112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13712 GND A2 word288 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13713 a_1106_n61686# a_1056_n66# a_974_n61686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13714 a_1106_n70064# a_1056_n66# a_842_n70064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13715 word790 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13716 a_1238_n120190# A5 a_842_n120190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13717 GND A4 word719 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13718 a_50_n84406# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13719 word406 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13720 a_2294_n7016# A1 a_2030_n7016# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13721 a_974_n92926# A6 a_578_n92926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13722 word435 a_2376_n66# a_2162_n61970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13723 GND A7 word290 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13724 GND A2 word817 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13725 a_50_n110960# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13726 a_1502_n137798# A4 a_1238_n137798# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13727 a_1370_n48480# a_1320_n66# a_1238_n48480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13728 GND A7 word620 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13729 a_842_n71342# a_792_n66# a_578_n71342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13730 a_974_n78442# A6 a_710_n78442# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13731 a_578_n22210# a_528_n66# a_446_n22210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13732 word333 a_2376_n66# a_2294_n47486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13733 a_1766_n96050# A3 a_1502_n96050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13734 word125 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13735 word184 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13736 a_182_n52314# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13737 a_314_n59414# a_264_n66# a_182_n59414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13738 GND A0 word252 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13739 GND A1 word269 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13740 a_182_n43936# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13741 word462 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13742 a_578_n91506# a_528_n66# a_446_n91506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13743 word1022 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13744 word963 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13745 a_1898_n73614# a_1848_n66# a_1766_n73614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13746 a_578_n30162# a_528_n66# a_446_n30162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13747 a_182_n29452# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13748 a_578_n21784# a_528_n66# a_446_n21784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13749 a_1238_n11702# A5 a_842_n11702# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13750 a_842_n101872# a_792_n66# a_578_n101872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13751 a_842_n31440# a_792_n66# a_578_n31440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13752 a_974_n38540# A6 a_710_n38540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13753 word895 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13754 word25 a_2376_n66# a_2294_n3750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13755 a_974_n60976# A6 a_578_n60976# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13756 GND A6 word516 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13757 word674 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13758 word760 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13759 a_50_n99316# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13760 a_578_n68644# a_528_n66# a_314_n68644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13761 GND A4 word455 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13762 a_314_n50326# a_264_n66# a_182_n50326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13763 word669 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13764 a_314_n41948# a_264_n66# a_182_n41948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13765 word599 a_2376_n66# a_2162_n85258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13766 a_50_n134248# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13767 a_50_n125870# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13768 a_1766_n64100# A3 a_1502_n64100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13769 GND A0 word518 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13770 a_1502_n63816# A4 a_1238_n63816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13771 word443 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13772 word816 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13773 word46 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13774 word384 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13775 word757 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13776 a_182_n11986# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13777 a_182_n20364# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13778 a_842_n86252# a_792_n66# a_710_n86252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13779 a_1898_n19228# a_1848_n66# a_1766_n19228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13780 word237 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13781 a_842_n108830# a_792_n66# a_578_n108830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13782 a_1898_n41664# a_1848_n66# a_1766_n41664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13783 a_1898_n50042# a_1848_n66# a_1634_n50042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13784 GND A0 word416 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13785 word506 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13786 word738 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13787 a_182_n58846# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13788 a_182_n67224# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13789 a_50_n81850# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13790 a_50_n90228# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13791 GND A3 word193 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13792 word447 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13793 word742 A0 a_2162_n105564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13794 GND A2 word600 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13795 a_1898_n88524# a_1848_n66# a_1634_n88524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13796 GND A2 word858 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13797 GND A5 word131 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13798 GND A6 word133 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13799 word727 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13800 GND A4 word289 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13801 GND A4 word230 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13802 a_1238_n1620# A5 a_974_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13803 a_842_n46350# a_792_n66# a_710_n46350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13804 word501 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13805 word860 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13806 a_1898_n10140# a_1848_n66# a_1766_n10140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13807 a_1634_n65804# a_1584_n66# a_1502_n65804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13808 a_974_n75886# A6 a_710_n75886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13809 a_182_n9146# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13810 a_50_n102298# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13811 GND A0 word352 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13812 word1023 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13813 a_314_n56858# a_264_n66# a_182_n56858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13814 a_314_n65236# a_264_n66# a_182_n65236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13815 a_1106_n123314# a_1056_n66# a_842_n123314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13816 a_1634_n115504# a_1584_n66# a_1502_n115504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13817 GND A4 word128 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13818 a_314_n111528# a_264_n66# a_50_n111528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13819 word503 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13820 a_1106_n114936# a_1056_n66# a_974_n114936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13821 GND A0 word682 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13822 a_2030_n7158# A2 a_1766_n7158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13823 word117 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13824 a_1502_n87104# A4 a_1106_n87104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13825 word1008 A0 a_2294_n143336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13826 word916 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13827 a_1502_n78726# A4 a_1106_n78726# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13828 a_182_n35274# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13829 GND A4 word616 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13830 word489 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13831 a_182_n26896# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13832 word220 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13833 word401 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13834 word993 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13835 word934 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13836 word902 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13837 a_1898_n56574# a_1848_n66# a_1634_n56574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13838 a_710_n7300# A7 a_446_n7300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13839 a_50_n96760# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13840 GND A3 word38 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13841 a_842_n14400# a_792_n66# a_710_n14400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13842 a_50_n140070# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13843 word241 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13844 a_974_n111954# A6 a_710_n111954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13845 word832 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13846 GND A2 word904 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13847 a_1634_n42232# a_1584_n66# a_1502_n42232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13848 word381 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13849 word613 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13850 word773 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13851 a_1634_n33854# a_1584_n66# a_1502_n33854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13852 GND A4 word335 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13853 GND A4 word394 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13854 word554 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13855 word425 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13856 word606 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13857 a_974_n99174# A6 a_578_n99174# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13858 word965 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13859 a_842_n123030# a_792_n66# a_710_n123030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13860 GND A6 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13861 a_1898_n25050# a_1848_n66# a_1634_n25050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13862 a_842_n83696# a_792_n66# a_710_n83696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13863 a_182_n64668# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13864 a_1502_n46776# A4 a_1238_n46776# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13865 a_1502_n55154# A4 a_1238_n55154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13866 a_314_n126438# a_264_n66# a_50_n126438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13867 word323 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13868 word264 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13869 GND A0 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13870 word446 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13871 a_1898_n94346# a_1848_n66# a_1766_n94346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13872 a_2030_n200# A2 a_1766_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13873 a_1502_n6448# A4 a_1106_n6448# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13874 word176 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13875 a_1898_n85968# a_1848_n66# a_1634_n85968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13876 word1021 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13877 word709 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13878 a_50_n73188# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13879 word325 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13880 word448 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13881 a_182_n6590# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13882 a_314_n62680# a_264_n66# a_182_n62680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13883 a_314_n71058# a_264_n66# a_182_n71058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13884 word97 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13885 GND A3 word561 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13886 GND A4 word169 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13887 word346 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13888 a_974_n135242# A6 a_578_n135242# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13889 a_1634_n112948# a_1584_n66# a_1370_n112948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13890 word740 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13891 GND A0 word664 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13892 word990 A0 a_2162_n140780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13893 GND A6 word779 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13894 a_1766_n121610# A3 a_1370_n121610# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13895 a_182_n41096# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13896 a_314_n48196# a_264_n66# a_182_n48196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13897 a_1106_n106274# a_1056_n66# a_842_n106274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13898 a_1370_n7158# a_1320_n66# a_1106_n7158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13899 GND A3 word339 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13900 a_1898_n62396# a_1848_n66# a_1766_n62396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13901 a_1766_n107126# A3 a_1370_n107126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13902 GND A9 word431 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13903 word888 A0 a_2294_n126296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13904 GND A3 word497 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13905 word551 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13906 GND A0 word52 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13907 word100 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13908 a_1634_n17240# a_1584_n66# a_1370_n17240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13909 a_2030_n17524# A2 a_1634_n17524# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13910 word205 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13911 word223 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13912 word873 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13913 GND A2 word945 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13914 GND A5 word277 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13915 word363 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13916 word814 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13917 word654 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13918 a_1238_n47344# A5 a_842_n47344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13919 word595 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13920 a_50_n88098# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13921 a_1238_n38966# A5 a_974_n38966# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13922 word612 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13923 word647 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13924 word693 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13925 word121 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13926 word424 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13927 word588 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13928 word261 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13929 word334 A0 a_2162_n47628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13930 a_182_n70490# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13931 a_314_n132260# a_264_n66# a_50_n132260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13932 word743 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13933 a_1106_n144046# a_1056_n66# a_842_n144046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13934 a_1634_n136236# a_1584_n66# a_1370_n136236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13935 a_1106_n135668# a_1056_n66# a_974_n135668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13936 word270 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13937 a_2162_n77732# a_2112_n66# a_2030_n77732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13938 word649 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13939 GND A5 word213 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13940 a_1898_n91790# a_1848_n66# a_1766_n91790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13941 GND A6 word943 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13942 GND A7 word796 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13943 a_1766_n136520# A3 a_1502_n136520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13944 GND A3 word114 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13945 a_2030_n124024# A2 a_1634_n124024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13946 a_2030_n46918# A2 a_1634_n46918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13947 a_314_n109398# a_264_n66# a_50_n109398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13948 GND A5 word543 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13949 word488 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13950 word326 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13951 a_578_n95198# a_528_n66# a_446_n95198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13952 a_1238_n85116# A5 a_842_n85116# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13953 a_1238_n76738# A5 a_974_n76738# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13954 GND A3 word661 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13955 GND A9 word477 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13956 a_2294_n75744# A1 a_1898_n75744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13957 GND A1 word801 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13958 word328 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13959 word527 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13960 word978 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13961 a_974_n132686# A6 a_578_n132686# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13962 a_1634_n54586# a_1584_n66# a_1370_n54586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13963 word700 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13964 word168 A0 a_2294_n24056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13965 a_2162_n108546# a_2112_n66# a_2030_n108546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13966 word1001 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13967 a_446_n27606# A8 a_182_n27606# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13968 a_1634_n104286# a_1584_n66# a_1370_n104286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13969 a_1370_n111812# a_1320_n66# a_1238_n111812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13970 GND A9 word255 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13971 word656 A0 a_2294_n93352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13972 word695 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13973 a_710_n41238# A7 a_314_n41238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13974 a_2030_n23346# A2 a_1766_n23346# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13975 a_446_n96902# A8 a_50_n96902# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13976 a_2030_n14968# A2 a_1634_n14968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13977 word281 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13978 word1005 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13979 word720 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13980 word222 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13981 GND A5 word259 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13982 GND A7 word842 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13983 word594 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13984 GND A3 word1012 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13985 GND A9 word311 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13986 a_1238_n140922# A5 a_842_n140922# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13987 a_2162_n14258# a_2112_n66# a_2030_n14258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13988 a_710_n79720# A7 a_446_n79720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13989 a_1634_n92358# a_1584_n66# a_1502_n92358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13990 GND A9 word252 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13991 GND A6 word24 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13992 a_1634_n83980# a_1584_n66# a_1502_n83980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13993 a_2030_n92642# A2 a_1634_n92642# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X13994 a_2162_n137940# a_2112_n66# a_2030_n137940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13995 word903 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13996 a_2294_n99032# A1 a_2030_n99032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13997 GND A8 word712 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X13998 a_1106_n141490# a_1056_n66# a_842_n141490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X13999 GND A8 word151 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14000 a_2162_n83554# a_2112_n66# a_2030_n83554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14001 a_1634_n133680# a_1584_n66# a_1502_n133680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14002 a_1898_n121184# a_1848_n66# a_1766_n121184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14003 word43 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14004 a_2294_n103718# A1 a_2030_n103718# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14005 word304 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14006 a_1634_n69496# a_1584_n66# a_1502_n69496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14007 a_710_n87672# A7 a_446_n87672# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14008 GND A6 word925 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14009 word245 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14010 GND A7 word778 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14011 a_1370_n126722# a_1320_n66# a_1106_n126722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14012 a_2294_n12270# A1 a_1898_n12270# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14013 GND A2 word153 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14014 a_2030_n52740# A2 a_1766_n52740# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14015 GND A5 word584 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14016 GND A5 word525 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14017 GND A3 word485 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14018 a_1238_n82560# A5 a_842_n82560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14019 GND A6 word823 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14020 word702 A0 a_2162_n99884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14021 a_2294_n81566# A1 a_1898_n81566# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14022 a_710_n47770# A7 a_314_n47770# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14023 GND A8 word39 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14024 word369 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14025 GND A3 word787 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14026 a_2030_n29878# A2 a_1766_n29878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14027 a_2030_n60692# A2 a_1634_n60692# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14028 word509 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14029 word787 a_2376_n66# a_2162_n111954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14030 a_1238_n68076# A5 a_842_n68076# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14031 word150 A0 a_2162_n21500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14032 GND A7 word112 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14033 GND A9 word416 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14034 a_446_n33428# A8 a_182_n33428# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14035 GND A1 word193 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14036 word570 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14037 GND A9 word27 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14038 word480 A0 a_2294_n68360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14039 word638 A0 a_2162_n90796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14040 word889 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14041 GND A8 word758 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14042 a_1898_n136094# a_1848_n66# a_1634_n136094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14043 a_2294_n127006# A1 a_1898_n127006# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14044 word746 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14045 a_1766_n84832# A3 a_1370_n84832# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14046 GND A1 word681 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14047 word105 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14048 a_2030_n20790# A2 a_1766_n20790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14049 a_842_n9998# a_792_n66# a_710_n9998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14050 GND A7 word58 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14051 GND A7 word883 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14052 GND A9 word135 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14053 GND A2 word258 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14054 word635 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14055 GND A9 word352 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14056 a_578_n138224# a_528_n66# a_314_n138224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14057 GND A4 word748 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14058 word42 A0 a_2162_n6164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14059 a_2030_n67650# A2 a_1634_n67650# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14060 a_578_n129846# a_528_n66# a_314_n129846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14061 a_446_n79862# A8 a_50_n79862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14062 GND A5 word981 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14063 word944 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14064 word91 a_2376_n66# a_2162_n13122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14065 a_1766_n53308# A3 a_1370_n53308# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14066 GND A3 word951 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14067 word951 a_2376_n66# a_2162_n135242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14068 word25 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14069 GND A8 word522 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14070 word856 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14071 word953 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14072 word675 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14073 GND A1 word456 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14074 a_974_n6874# A6 a_710_n6874# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14075 a_1766_n52882# A3 a_1370_n52882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14076 GND A5 word917 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14077 GND A1 word725 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14078 a_1502_n141206# A4 a_1106_n141206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14079 a_1502_n132828# A4 a_1106_n132828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14080 a_1106_n33854# a_1056_n66# a_842_n33854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14081 a_1106_n42232# a_1056_n66# a_974_n42232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14082 a_578_n25902# a_528_n66# a_446_n25902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14083 a_1370_n43510# a_1320_n66# a_1106_n43510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14084 a_578_n106274# a_528_n66# a_446_n106274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14085 a_2030_n35700# A2 a_1634_n35700# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14086 GND A5 word464 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14087 a_1238_n139218# A5 a_842_n139218# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14088 GND A7 word94 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14089 word719 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14090 GND A9 word457 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14091 a_1502_n118344# A4 a_1238_n118344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14092 GND A3 word726 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14093 a_1502_n109966# A4 a_1238_n109966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14094 a_1766_n21358# A3 a_1370_n21358# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14095 word698 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14096 GND A9 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14097 GND A0 word834 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14098 word207 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14099 a_446_n86110# A8 a_50_n86110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14100 word137 a_2376_n66# a_2294_n19654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14101 a_1766_n59840# A3 a_1502_n59840# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14102 GND A8 word238 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14103 word728 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14104 GND A7 word582 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14105 a_1238_n138792# A5 a_842_n138792# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14106 a_446_n16388# A8 a_182_n16388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14107 word146 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14108 a_1370_n89944# a_1320_n66# a_1106_n89944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14109 a_1370_n98322# a_1320_n66# a_1106_n98322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14110 GND A7 word40 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14111 a_1106_n80004# a_1056_n66# a_974_n80004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14112 word860 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14113 GND A8 word627 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14114 a_1238_n130130# A5 a_974_n130130# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14115 GND A2 word299 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14116 a_1106_n71626# a_1056_n66# a_842_n71626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14117 a_2030_n142200# A2 a_1634_n142200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14118 word769 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14119 a_578_n144046# a_528_n66# a_314_n144046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14120 a_1502_n100878# A4 a_1238_n100878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14121 a_578_n135668# a_528_n66# a_314_n135668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14122 word58 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14123 a_446_n85684# A8 a_50_n85684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14124 a_446_n94062# A8 a_50_n94062# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14125 GND A1 word561 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14126 word634 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14127 a_1370_n11560# a_1320_n66# a_1238_n11560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14128 word575 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14129 GND A5 word963 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14130 word985 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14131 a_974_n41522# A6 a_710_n41522# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14132 word505 a_2376_n66# a_2294_n71910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14133 GND A7 word360 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14134 word73 a_2376_n66# a_2294_n10566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14135 word916 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14136 GND A3 word992 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14137 GND A1 word988 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14138 GND A3 word933 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14139 GND A2 word138 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14140 a_1370_n58420# a_1320_n66# a_1238_n58420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14141 word857 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14142 word473 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14143 a_2162_n135100# a_2112_n66# a_1898_n135100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14144 word933 a_2376_n66# a_2294_n132686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14145 word403 a_2376_n66# a_2162_n57426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14146 word414 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14147 a_1370_n80856# a_1320_n66# a_1106_n80856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14148 GND A8 word563 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14149 a_50_n106416# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14150 a_1634_n6732# a_1584_n66# a_1502_n6732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14151 GND A0 word322 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14152 a_1766_n27890# A3 a_1502_n27890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14153 GND A1 word280 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14154 GND A1 word497 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14155 GND A7 word357 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14156 a_1370_n66372# a_1320_n66# a_1238_n66372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14157 a_1106_n17240# a_1056_n66# a_842_n17240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14158 a_1370_n57994# a_1320_n66# a_1238_n57994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14159 a_2294_n139360# A1 a_1898_n139360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14160 a_578_n31724# a_528_n66# a_446_n31724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14161 GND A1 word64 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14162 word251 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14163 a_1106_n86536# a_1056_n66# a_842_n86536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14164 word965 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14165 GND A5 word797 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14166 a_1502_n124166# A4 a_1106_n124166# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14167 GND A4 word835 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14168 a_1106_n25192# a_1056_n66# a_974_n25192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14169 a_710_n112380# A7 a_314_n112380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14170 a_1502_n115788# A4 a_1106_n115788# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14171 GND A3 word67 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14172 word680 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14173 a_1370_n26470# a_1320_n66# a_1106_n26470# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14174 a_50_n135810# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14175 a_974_n56432# A6 a_578_n56432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14176 GND A1 word605 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14177 word1021 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14178 word886 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14179 GND A0 word156 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14180 word827 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14181 a_182_n30304# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14182 a_314_n37404# a_264_n66# a_182_n37404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14183 GND A6 word50 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14184 GND A4 word581 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14185 GND A8 word668 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14186 a_182_n21926# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14187 GND A6 word305 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14188 a_842_n87814# a_792_n66# a_710_n87814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14189 GND A8 word609 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14190 GND A0 word486 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14191 a_1370_n144898# a_1320_n66# a_1106_n144898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14192 word867 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14193 a_578_n141490# a_528_n66# a_314_n141490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14194 a_710_n2330# A7 a_446_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14195 GND A1 word661 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14196 GND A7 word521 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14197 word812 A0 a_2294_n115504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14198 a_50_n143762# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14199 a_2030_n1762# A2 a_1634_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14200 a_1238_n113090# A5 a_974_n113090# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14201 a_578_n55012# a_528_n66# a_314_n55012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14202 a_1106_n54586# a_1056_n66# a_842_n54586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14203 a_842_n126722# a_792_n66# a_710_n126722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14204 a_50_n77306# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14205 a_974_n94204# A6 a_578_n94204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14206 GND A5 word902 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14207 GND A6 word691 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14208 a_50_n112238# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14209 word385 a_2376_n66# a_2294_n54870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14210 GND A0 word422 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14211 a_710_n127290# A7 a_314_n127290# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14212 a_50_n103860# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14213 a_974_n24482# A6 a_578_n24482# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14214 a_1766_n42090# A3 a_1502_n42090# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14215 GND A1 word380 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14216 GND A4 word139 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14217 GND A4 word198 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14218 a_1502_n41806# A4 a_1106_n41806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14219 GND A0 word980 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14220 GND A4 word356 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14221 a_1370_n72194# a_1320_n66# a_1106_n72194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14222 a_842_n64242# a_792_n66# a_578_n64242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14223 word141 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14224 word927 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14225 GND A0 word202 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14226 word351 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14227 GND A4 word686 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14228 a_182_n36836# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14229 a_182_n45214# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14230 a_1502_n18944# A4 a_1238_n18944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14231 GND A6 word410 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14232 word412 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14233 GND A6 word568 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14234 GND A7 word626 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14235 a_182_n1620# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14236 word766 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14237 a_578_n23062# a_528_n66# a_446_n23062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14238 GND A4 word75 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14239 a_974_n62254# A6 a_578_n62254# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14240 word843 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14241 word219 a_2376_n66# a_2162_n31298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14242 word287 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14243 a_1106_n69496# a_1056_n66# a_842_n69496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14244 word624 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14245 GND A6 word407 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14246 word868 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14247 a_314_n43226# a_264_n66# a_182_n43226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14248 word619 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14249 GND A4 word37 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14250 word549 a_2376_n66# a_2294_n78158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14251 GND A8 word650 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14252 a_50_n127148# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14253 a_974_n39392# A6 a_710_n39392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14254 GND A7 word345 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14255 a_50_n118770# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14256 a_842_n32292# a_792_n66# a_578_n32292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14257 GND A0 word468 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14258 GND A1 word485 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14259 a_1766_n3182# A3 a_1370_n3182# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14260 a_1502_n56716# A4 a_1238_n56716# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14261 word393 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14262 word794 A0 a_2162_n112948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14263 a_182_n13264# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14264 GND A4 word461 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14265 word334 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14266 GND A6 word185 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14267 word246 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14268 word779 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14269 word187 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14270 word747 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14271 a_50_n83128# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14272 a_50_n74750# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14273 a_314_n135952# a_264_n66# a_50_n135952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14274 a_974_n91648# A6 a_578_n91648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14275 a_1106_n98890# a_1056_n66# a_974_n98890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14276 word86 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14277 a_578_n99316# a_528_n66# a_446_n99316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14278 GND A6 word673 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14279 a_314_n72620# a_264_n66# a_182_n72620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14280 a_1634_n20222# a_1584_n66# a_1502_n20222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14281 word167 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14282 a_578_n29594# a_528_n66# a_446_n29594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14283 a_1238_n19512# A5 a_974_n19512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14284 GND A4 word239 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14285 GND A3 word631 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14286 word42 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14287 a_842_n70064# a_792_n66# a_578_n70064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14288 a_1634_n58704# a_1584_n66# a_1370_n58704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14289 a_974_n77164# A6 a_710_n77164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14290 a_842_n101020# a_792_n66# a_578_n101020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14291 a_314_n58136# a_264_n66# a_182_n58136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14292 GND A0 word302 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14293 a_182_n42658# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14294 a_314_n49758# a_264_n66# a_182_n49758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14295 a_182_n51036# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14296 GND A2 word32 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14297 a_1502_n24766# A4 a_1106_n24766# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14298 a_1502_n33144# A4 a_1106_n33144# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14299 a_1106_n107836# a_1056_n66# a_842_n107836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14300 a_1634_n108404# a_1584_n66# a_1370_n108404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14301 a_1106_n116214# a_1056_n66# a_974_n116214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14302 word453 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14303 a_1370_n8720# a_1320_n66# a_1106_n8720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14304 word291 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14305 a_1898_n72336# a_1848_n66# a_1634_n72336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14306 word954 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14307 a_1238_n2472# A5 a_974_n2472# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14308 word604 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14309 word663 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14310 word958 A0 a_2162_n136236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14311 word807 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14312 a_1238_n10424# A5 a_842_n10424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14313 GND A3 word567 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14314 a_842_n100594# a_792_n66# a_578_n100594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14315 a_182_n28174# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14316 word943 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14317 a_182_n19796# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14318 word884 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14319 a_578_n67366# a_528_n66# a_314_n67366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14320 word665 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14321 a_50_n98038# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14322 word74 A0 a_2162_n10708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14323 a_578_n58988# a_528_n66# a_314_n58988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14324 a_1238_n48906# A5 a_842_n48906# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14325 a_314_n40670# a_264_n66# a_182_n40670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14326 a_50_n89660# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14327 word57 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14328 GND A3 word406 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14329 a_2294_n47912# A1 a_2030_n47912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14330 a_974_n113232# A6 a_710_n113232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14331 a_2162_n40812# a_2112_n66# a_1898_n40812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14332 word331 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14333 a_1634_n26754# a_1584_n66# a_1370_n26754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14334 word375 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14335 word498 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14336 word556 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14337 word660 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14338 a_1898_n116924# a_1848_n66# a_1766_n116924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14339 a_1238_n9430# A5 a_842_n9430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14340 word228 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14341 word438 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14342 a_182_n57568# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14343 a_314_n119338# a_264_n66# a_50_n119338# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14344 a_314_n141774# a_264_n66# a_50_n141774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14345 a_710_n13406# A7 a_446_n13406# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14346 a_578_n96760# a_528_n66# a_446_n96760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14347 a_1898_n87246# a_1848_n66# a_1766_n87246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14348 word718 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14349 GND A3 word672 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14350 word492 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14351 a_710_n82702# A7 a_446_n82702# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14352 word1014 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14353 word1012 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14354 a_2162_n140922# a_2112_n66# a_1898_n140922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14355 a_314_n55580# a_264_n66# a_182_n55580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14356 a_314_n110250# a_264_n66# a_50_n110250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14357 a_1634_n105848# a_1584_n66# a_1502_n105848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14358 word115 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14359 a_2162_n55722# a_2112_n66# a_1898_n55722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14360 word435 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14361 word494 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14362 a_974_n128142# A6 a_578_n128142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14363 GND A0 word614 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14364 word995 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14365 word108 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14366 a_1502_n77448# A4 a_1106_n77448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14367 word940 A0 a_2294_n133680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14368 word662 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14369 word480 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14370 a_1766_n114510# A3 a_1502_n114510# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14371 word603 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14372 word925 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14373 word171 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14374 GND A5 word329 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14375 a_1898_n55296# a_1848_n66# a_1766_n55296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14376 a_1238_n54728# A5 a_974_n54728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14377 GND A9 word381 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14378 a_842_n144898# a_792_n66# a_578_n144898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14379 word838 A0 a_2162_n119196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14380 GND A9 word322 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14381 a_2162_n15820# a_2112_n66# a_1898_n15820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14382 a_2294_n53734# A1 a_2030_n53734# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14383 word232 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14384 a_2294_n62112# A1 a_1898_n62112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14385 a_974_n110676# A6 a_710_n110676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14386 word823 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14387 word764 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14388 a_710_n50752# A7 a_314_n50752# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14389 word313 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14390 word545 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14391 word846 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14392 word19 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14393 a_1898_n122746# a_1848_n66# a_1634_n122746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14394 word374 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14395 a_1634_n79436# a_1584_n66# a_1502_n79436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14396 a_2162_n23772# a_2112_n66# a_1898_n23772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14397 word315 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14398 a_1634_n18092# a_1584_n66# a_1370_n18092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14399 GND A3 word225 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14400 GND A7 word848 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14401 a_1634_n129136# a_1584_n66# a_1502_n129136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14402 a_182_n63390# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14403 word442 A0 a_2162_n62964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14404 a_314_n125160# a_264_n66# a_50_n125160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14405 word7 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14406 a_1502_n5170# A4 a_1106_n5170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14407 word378 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14408 a_1898_n93068# a_1848_n66# a_1634_n93068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14409 a_710_n10850# A7 a_446_n10850# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14410 a_1238_n31156# A5 a_842_n31156# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14411 word371 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14412 a_1238_n22778# A5 a_974_n22778# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14413 a_2030_n108546# A2 a_1634_n108546# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14414 GND A9 word156 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14415 a_1634_n70348# a_1584_n66# a_1502_n70348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14416 word579 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14417 GND A9 word97 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14418 a_2294_n21784# A1 a_2030_n21784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14419 a_2030_n70632# A2 a_1766_n70632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14420 GND A5 word651 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14421 a_2030_n130982# A2 a_1634_n130982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14422 a_2162_n124308# a_2112_n66# a_2030_n124308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14423 a_2162_n115930# a_2112_n66# a_1898_n115930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14424 word701 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14425 word147 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14426 word220 A0 a_2294_n31440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14427 word748 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14428 GND A9 word486 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14429 a_2162_n39108# a_2112_n66# a_2030_n39108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14430 a_2294_n77022# A1 a_1898_n77022# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14431 a_1634_n120048# a_1584_n66# a_1502_n120048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14432 word337 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14433 a_1766_n137372# A3 a_1502_n137372# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14434 a_974_n1904# A6 a_710_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14435 a_1634_n47486# a_1584_n66# a_1502_n47486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14436 a_1502_n83270# A4 a_1238_n83270# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14437 word892 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14438 a_578_n101304# a_528_n66# a_446_n101304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14439 a_2162_n123882# a_2112_n66# a_1898_n123882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14440 word420 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14441 a_2162_n38682# a_2112_n66# a_1898_n38682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14442 word637 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14443 word606 A0 a_2162_n86252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14444 GND A9 word422 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14445 GND A9 word205 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14446 a_2162_n30020# a_2112_n66# a_2030_n30020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14447 a_2294_n37120# A1 a_1898_n37120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14448 GND A9 word363 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14449 a_2030_n137940# A2 a_1634_n137940# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14450 a_446_n89802# A8 a_50_n89802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14451 word483 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14452 word542 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14453 a_2030_n16246# A2 a_1766_n16246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14454 word214 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14455 a_1898_n99600# a_1848_n66# a_1634_n99600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14456 GND A5 word209 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14457 GND A5 word268 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14458 word955 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14459 word172 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14460 a_1238_n37688# A5 a_974_n37688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14461 a_1238_n46066# A5 a_842_n46066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14462 GND A1 word1017 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14463 VDD A6 a_792_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X14464 a_2162_n90938# a_2112_n66# a_1898_n90938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14465 GND A9 word261 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14466 GND A9 word202 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14467 GND A3 word962 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14468 a_446_n11418# A8 a_182_n11418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14469 a_2294_n45072# A1 a_1898_n45072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14470 a_2030_n85542# A2 a_1634_n85542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14471 word625 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14472 a_2162_n139218# a_2112_n66# a_2030_n139218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14473 a_2294_n36694# A1 a_2030_n36694# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14474 a_1634_n76880# a_1584_n66# a_1370_n76880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14475 word1011 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14476 word640 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14477 a_1106_n134390# a_1056_n66# a_974_n134390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14478 word726 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14479 a_1634_n126580# a_1584_n66# a_1370_n126580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14480 GND A8 word101 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14481 a_446_n107552# A8 a_50_n107552# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14482 a_446_n80714# A8 a_50_n80714# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14483 GND A5 word145 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14484 word254 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14485 a_446_n10992# A8 a_182_n10992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14486 GND A2 word162 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14487 a_2030_n54018# A2 a_1634_n54018# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14488 a_578_n107836# a_528_n66# a_446_n107836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14489 a_2030_n45640# A2 a_1766_n45640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14490 GND A5 word475 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14491 GND A5 word534 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14492 a_2030_n105990# A2 a_1634_n105990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14493 a_2162_n130130# a_2112_n66# a_2030_n130130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14494 a_1238_n75460# A5 a_974_n75460# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14495 word730 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14496 GND A9 word468 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14497 a_1502_n119906# A4 a_1238_n119906# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14498 a_1766_n22920# A3 a_1502_n22920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14499 a_710_n49048# A7 a_314_n49048# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14500 GND A8 word48 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14501 GND A3 word737 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14502 GND A1 word792 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14503 word459 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14504 a_1238_n101872# A5 a_842_n101872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14505 word737 a_2376_n66# a_2294_n104854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14506 a_2030_n53592# A2 a_1634_n53592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14507 a_2162_n107268# a_2112_n66# a_2030_n107268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14508 word992 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14509 word100 A0 a_2294_n14400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14510 a_710_n626# A7 a_446_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14511 word798 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14512 a_446_n26328# A8 a_182_n26328# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14513 a_446_n17950# A8 a_182_n17950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14514 GND A1 word29 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14515 GND A1 word301 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14516 GND A8 word767 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14517 word839 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14518 GND A8 word206 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14519 word588 A0 a_2294_n83696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14520 a_1502_n110818# A4 a_1238_n110818# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14521 a_446_n95624# A8 a_50_n95624# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14522 word997 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14523 a_2030_n22068# A2 a_1634_n22068# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14524 a_1766_n77732# A3 a_1502_n77732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14525 a_2294_n142342# A1 a_2030_n142342# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14526 GND A2 word267 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14527 GND A7 word833 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14528 word986 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14529 word143 a_2376_n66# a_2162_n20506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14530 GND A2 word208 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14531 word585 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14532 word927 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14533 GND A9 word302 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14534 a_1106_n7868# a_1056_n66# a_974_n7868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14535 a_2030_n91364# A2 a_1766_n91364# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14536 word1003 a_2376_n66# a_2162_n142626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14537 a_710_n17098# A7 a_446_n17098# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14538 GND A6 word15 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14539 word543 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14540 GND A8 word574 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14541 a_1766_n46208# A3 a_1502_n46208# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14542 GND A8 word142 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14543 GND A8 word703 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14544 word1005 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14545 GND A3 word901 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14546 word775 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14547 GND A8 word83 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14548 a_2162_n73898# a_2112_n66# a_1898_n73898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14549 a_2162_n82276# a_2112_n66# a_2030_n82276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14550 a_2294_n89376# A1 a_1898_n89376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14551 a_2294_n102440# A1 a_2030_n102440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14552 word901 a_2376_n66# a_2294_n128142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14553 GND A1 word897 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14554 a_1370_n76312# a_1320_n66# a_1238_n76312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14555 a_710_n86394# A7 a_446_n86394# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14556 a_446_n104996# A8 a_50_n104996# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14557 word295 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14558 a_1370_n67934# a_1320_n66# a_1238_n67934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14559 GND A1 word76 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14560 GND A2 word144 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14561 a_1370_n125444# a_1320_n66# a_1106_n125444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14562 GND A7 word266 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14563 a_974_n8152# A6 a_710_n8152# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14564 a_1766_n45782# A3 a_1502_n45782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14565 a_2294_n110392# A1 a_2030_n110392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14566 GND A2 word474 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14567 a_1502_n134106# A4 a_1106_n134106# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14568 GND A4 word905 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14569 a_1106_n35132# a_1056_n66# a_842_n35132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14570 GND A9 word509 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14571 a_710_n122320# A7 a_314_n122320# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14572 a_1106_n26754# a_1056_n66# a_974_n26754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14573 GND A8 word30 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14574 a_2294_n80288# A1 a_1898_n80288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14575 a_578_n18802# a_528_n66# a_446_n18802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14576 a_2030_n28600# A2 a_1634_n28600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14577 a_1370_n36410# a_1320_n66# a_1106_n36410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14578 word318 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14579 a_2162_n113090# a_2112_n66# a_2030_n113090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14580 word780 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14581 a_446_n32150# A8 a_182_n32150# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14582 a_1766_n14258# A3 a_1502_n14258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14583 GND A1 word125 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14584 GND A1 word184 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14585 a_2030_n97896# A2 a_1766_n97896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14586 GND A4 word961 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14587 GND A8 word679 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14588 a_710_n121894# A7 a_314_n121894# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14589 a_1370_n44362# a_1320_n66# a_1106_n44362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14590 a_1370_n35984# a_1320_n66# a_1106_n35984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14591 a_446_n79010# A8 a_50_n79010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14592 GND A8 word247 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14593 a_2162_n97186# a_2112_n66# a_2030_n97186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14594 GND A7 word532 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14595 GND A7 word591 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14596 GND A8 word749 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14597 GND A0 word942 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14598 GND A8 word188 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14599 GND A1 word672 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14600 a_2294_n117350# A1 a_2030_n117350# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14601 GND A7 word49 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14602 word810 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14603 GND A6 word431 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14604 GND A4 word739 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14605 GND A2 word249 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14606 a_1502_n102156# A4 a_1238_n102156# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14607 a_578_n128568# a_528_n66# a_314_n128568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14608 a_446_n7442# A8 a_182_n7442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14609 word584 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14610 a_446_n78584# A8 a_50_n78584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14611 word525 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14612 GND A5 word972 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14613 word455 a_2376_n66# a_2162_n64810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14614 GND A7 word310 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14615 GND A0 word720 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14616 GND A5 word913 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14617 a_2294_n95198# A1 a_1898_n95198# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14618 a_2162_n3466# a_2112_n66# a_1898_n3466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14619 word807 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14620 word866 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14621 GND A3 word883 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14622 word883 a_2376_n66# a_2162_n125586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14623 GND A8 word513 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14624 a_842_n65804# a_792_n66# a_578_n65804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14625 GND A7 word366 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14626 word511 a_2376_n66# a_2162_n72762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14627 a_1370_n131266# a_1320_n66# a_1238_n131266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14628 GND A0 word776 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14629 a_50_n121752# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14630 GND A0 word272 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14631 GND A7 word307 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14632 a_974_n5596# A6 a_710_n5596# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14633 GND A9 word64 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14634 GND A2 word515 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14635 GND A5 word849 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14636 a_578_n33002# a_528_n66# a_446_n33002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14637 a_1106_n32576# a_1056_n66# a_842_n32576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14638 a_842_n104712# a_792_n66# a_578_n104712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14639 a_1766_n98464# A3 a_1370_n98464# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14640 word836 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14641 a_578_n24624# a_528_n66# a_446_n24624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14642 word289 a_2376_n66# a_2294_n41238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14643 word300 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14644 a_1106_n79436# a_1056_n66# a_974_n79436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14645 GND A6 word536 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14646 GND A7 word85 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14647 GND A2 word571 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14648 a_1106_n18092# a_1056_n66# a_842_n18092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14649 GND A1 word225 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14650 GND A4 word1002 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14651 a_50_n128710# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14652 GND A7 word573 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14653 word971 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14654 a_1766_n4744# A3 a_1502_n4744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14655 a_842_n33854# a_792_n66# a_578_n33854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14656 word719 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14657 a_182_n23204# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14658 GND A0 word106 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14659 a_182_n14826# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14660 a_1106_n70348# a_1056_n66# a_842_n70348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14661 GND A8 word559 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14662 word952 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14663 GND A2 word290 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14664 a_1106_n61970# a_1056_n66# a_974_n61970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14665 word758 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14666 a_578_n134390# a_528_n66# a_314_n134390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14667 a_50_n136662# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14668 word467 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14669 word762 A0 a_2162_n108404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14670 a_446_n4886# A8 a_182_n4886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14671 word49 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14672 GND A1 word552 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14673 a_974_n40244# A6 a_710_n40244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14674 GND A6 word311 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14675 a_842_n119622# a_792_n66# a_710_n119622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14676 a_710_n3182# A7 a_446_n3182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14677 a_50_n92642# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14678 a_974_n78726# A6 a_710_n78726# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14679 a_842_n71626# a_792_n66# a_578_n71626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14680 word462 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14681 word985 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14682 a_50_n105138# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14683 word335 a_2376_n66# a_2162_n47770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14684 GND A0 word372 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14685 a_842_n10282# a_792_n66# a_710_n10282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14686 a_842_n48764# a_792_n66# a_710_n48764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14687 a_578_n30446# a_528_n66# a_446_n30446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14688 word877 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14689 a_182_n38114# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14690 a_1898_n12554# a_1848_n66# a_1766_n12554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14691 word242 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14692 a_182_n29736# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14693 GND A3 word146 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14694 GND A2 word395 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14695 a_314_n113942# a_264_n66# a_50_n113942# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14696 GND A5 word788 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14697 a_578_n68928# a_528_n66# a_314_n68928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14698 GND A6 word518 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14699 a_314_n50610# a_264_n66# a_182_n50610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14700 a_2030_n9572# A2 a_1766_n9572# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14701 a_842_n17240# a_792_n66# a_710_n17240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14702 word237 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14703 a_974_n55154# A6 a_578_n55154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14704 GND A6 word416 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14705 word169 a_2376_n66# a_2294_n24198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14706 GND A0 word88 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14707 word818 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14708 word759 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14709 a_182_n2472# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14710 a_182_n20648# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14711 a_1502_n11134# A4 a_1238_n11134# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14712 a_842_n86536# a_792_n66# a_710_n86536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14713 a_1370_n94488# a_1320_n66# a_1238_n94488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14714 GND A8 word600 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14715 word858 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14716 a_1898_n768# a_1848_n66# a_1766_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14717 GND A0 word418 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14718 word657 a_2376_n66# a_2294_n93494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14719 word799 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14720 a_182_n67508# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14721 a_50_n142484# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14722 a_1898_n41948# a_1848_n66# a_1766_n41948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14723 word508 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14724 word711 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14725 word744 A0 a_2294_n105848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14726 a_2294_n200# A1 a_2030_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14727 word36 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14728 GND A0 word576 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14729 word501 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14730 GND A6 word135 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14731 word137 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14732 word196 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14733 word729 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14734 word442 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14735 GND A9 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14736 word982 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14737 a_842_n125444# a_792_n66# a_710_n125444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14738 a_50_n76028# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14739 word347 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14740 a_2294_n25902# A1 a_1898_n25902# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14741 word503 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14742 a_314_n128852# a_264_n66# a_50_n128852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14743 GND A6 word682 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14744 a_182_n9430# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14745 word71 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14746 a_1634_n13122# a_1584_n66# a_1370_n13122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14747 GND A0 word354 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14748 a_314_n65520# a_264_n66# a_182_n65520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14749 word117 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14750 GND A2 word857 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14751 GND A4 word130 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14752 word566 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14753 GND A0 word684 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14754 word505 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14755 a_974_n129704# A6 a_578_n129704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14756 a_842_n54586# a_792_n66# a_710_n54586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14757 word342 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14758 word1010 A0 a_2162_n143620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14759 word918 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14760 a_1898_n1194# a_1848_n66# a_1766_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14761 GND A2 word41 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14762 word283 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14763 GND A4 word618 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14764 GND A4 word677 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14765 a_1106_n109114# a_1056_n66# a_842_n109114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14766 a_182_n35558# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14767 word403 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14768 a_1898_n56858# a_1848_n66# a_1634_n56858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14769 word908 A0 a_2294_n129136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14770 GND A3 word517 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14771 word757 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14772 a_1502_n86962# A4 a_1106_n86962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14773 a_1766_n132402# A3 a_1502_n132402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14774 word243 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14775 word893 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14776 a_1634_n42516# a_1584_n66# a_1502_n42516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14777 word615 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14778 word834 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14779 a_1106_n100026# a_1056_n66# a_974_n100026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14780 word800 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14781 a_974_n99458# A6 a_578_n99458# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14782 a_842_n83980# a_792_n66# a_710_n83980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14783 a_1634_n19654# a_1584_n66# a_1502_n19654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14784 a_1502_n55438# A4 a_1238_n55438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14785 GND A0 word400 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14786 word512 A0 a_2294_n72904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14787 word844 A0 a_2294_n120048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14788 GND A4 word452 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14789 word671 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14790 word325 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14791 a_1898_n118202# a_1848_n66# a_1634_n118202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14792 GND A0 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14793 a_1898_n109824# a_1848_n66# a_1766_n109824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14794 a_842_n69496# a_792_n66# a_578_n69496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14795 word178 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14796 word1023 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14797 word441 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14798 GND A3 word134 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14799 a_842_n122888# a_792_n66# a_710_n122888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14800 GND A3 word292 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14801 a_314_n143052# a_264_n66# a_50_n143052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14802 GND A9 word167 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14803 word77 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14804 a_2294_n40102# A1 a_2030_n40102# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14805 word346 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14806 a_1634_n71910# a_1584_n66# a_1370_n71910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14807 a_578_n98038# a_528_n66# a_446_n98038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14808 a_314_n134674# a_264_n66# a_50_n134674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14809 a_1766_n100452# A3 a_1502_n100452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14810 GND A6 word664 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14811 word217 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14812 word666 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14813 a_1634_n10566# a_1584_n66# a_1502_n10566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14814 word348 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14815 a_1898_n100736# a_1848_n66# a_1766_n100736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14816 a_1766_n138934# A3 a_1370_n138934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14817 a_974_n135526# A6 a_578_n135526# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14818 a_710_n75602# A7 a_446_n75602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14819 word383 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14820 a_1502_n93210# A4 a_1238_n93210# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14821 word160 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14822 word962 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14823 a_314_n48480# a_264_n66# a_182_n48480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14824 GND A3 word70 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14825 a_182_n41380# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14826 a_1502_n23488# A4 a_1106_n23488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14827 a_1106_n106558# a_1056_n66# a_842_n106558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14828 word444 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14829 word282 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14830 word385 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14831 word223 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14832 a_1238_n1194# A5 a_974_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14833 word595 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14834 a_1766_n107410# A3 a_1370_n107410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14835 word890 A0 a_2162_n126580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14836 GND A4 word557 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14837 a_1502_n92784# A4 a_1238_n92784# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14838 GND A0 word54 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14839 GND A5 word279 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14840 word875 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14841 a_578_n66088# a_528_n66# a_314_n66088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14842 a_1238_n47628# A5 a_842_n47628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14843 a_1238_n56006# A5 a_974_n56006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14844 word546 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14845 a_842_n137798# a_792_n66# a_578_n137798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14846 GND A9 word331 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14847 GND A9 word272 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14848 word123 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14849 word590 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14850 a_1766_n106984# A3 a_1370_n106984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14851 word263 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14852 GND A0 word500 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14853 a_710_n43652# A7 a_314_n43652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14854 a_1502_n61260# A4 a_1106_n61260# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14855 a_1106_n144330# a_1056_n66# a_842_n144330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14856 word737 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14857 a_1898_n115646# a_1848_n66# a_1634_n115646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14858 word219 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14859 word611 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14860 a_446_n20932# A8 a_182_n20932# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14861 GND A5 word215 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14862 a_1634_n94772# a_1584_n66# a_1370_n94772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14863 GND A7 word798 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14864 a_182_n56290# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14865 a_1502_n38398# A4 a_1238_n38398# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14866 a_314_n118060# a_264_n66# a_50_n118060# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14867 a_2030_n124308# A2 a_1634_n124308# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14868 a_2294_n15110# A1 a_2030_n15110# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14869 word392 A0 a_2294_n55864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14870 a_1634_n144472# a_1584_n66# a_1370_n144472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14871 word387 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14872 a_314_n140496# a_264_n66# a_50_n140496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14873 word490 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14874 word801 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14875 a_710_n12128# A7 a_446_n12128# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14876 word700 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14877 GND A3 word663 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14878 a_2294_n84406# A1 a_2030_n84406# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14879 GND A6 word942 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14880 word980 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14881 GND A9 word106 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14882 a_974_n132970# A6 a_578_n132970# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14883 a_1238_n111812# A5 a_974_n111812# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14884 a_2294_n23062# A1 a_2030_n23062# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14885 a_710_n81424# A7 a_446_n81424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14886 a_1634_n63248# a_1584_n66# a_1370_n63248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14887 word529 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14888 GND A5 word601 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14889 word1003 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14890 word170 A0 a_2162_n24340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14891 a_1238_n93352# A5 a_974_n93352# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14892 a_1238_n84974# A5 a_842_n84974# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14893 word695 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14894 a_1634_n104570# a_1584_n66# a_1370_n104570# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14895 a_2162_n54444# a_2112_n66# a_1898_n54444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14896 word99 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14897 word658 A0 a_2162_n93636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14898 word842 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14899 a_2030_n32008# A2 a_1766_n32008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14900 word226 A0 a_2162_n32292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14901 word594 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14902 a_2294_n143904# A1 a_1898_n143904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14903 GND A5 word320 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14904 a_446_n35842# A8 a_182_n35842# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14905 word556 A0 a_2294_n79152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14906 GND A9 word372 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14907 a_2030_n139218# A2 a_1766_n139218# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14908 word62 A0 a_2162_n9004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14909 GND A3 word438 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14910 GND A9 word313 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14911 GND A6 word776 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14912 a_2294_n52456# A1 a_2030_n52456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14913 a_1766_n121184# A3 a_1370_n121184# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14914 word905 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14915 word122 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14916 a_1634_n31298# a_1584_n66# a_1370_n31298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14917 word245 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14918 GND A8 word153 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14919 GND A8 word212 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14920 GND A3 word912 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14921 word836 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14922 a_1898_n121468# a_1848_n66# a_1766_n121468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14923 word365 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14924 a_1634_n69780# a_1584_n66# a_1502_n69780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14925 a_710_n87956# A7 a_446_n87956# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14926 a_2030_n138792# A2 a_1766_n138792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14927 word492 A0 a_2294_n70064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14928 GND A7 word780 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14929 word961 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14930 a_2030_n130130# A2 a_1766_n130130# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14931 a_1106_n127290# a_1056_n66# a_842_n127290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14932 a_2162_n69354# a_2112_n66# a_1898_n69354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14933 GND A7 word336 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14934 a_1634_n119480# a_1584_n66# a_1502_n119480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14935 a_446_n73614# A8 a_50_n73614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14936 a_1766_n55722# A3 a_1502_n55722# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14937 GND A5 word154 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14938 GND A6 word825 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14939 GND A5 word95 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14940 GND A2 word112 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14941 a_1238_n21500# A5 a_974_n21500# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14942 GND A7 word11 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14943 a_578_n109114# a_528_n66# a_446_n109114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14944 GND A3 word645 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14945 word699 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14946 GND A3 word848 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14947 a_2030_n107268# A2 a_1766_n107268# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14948 GND A9 word147 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14949 GND A9 word88 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14950 word692 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14951 word329 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14952 GND A5 word583 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14953 GND A5 word642 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14954 word739 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14955 GND A9 word418 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14956 a_2294_n67366# A1 a_2030_n67366# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14957 a_2162_n60266# a_2112_n66# a_1898_n60266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14958 GND A9 word29 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14959 a_1370_n54302# a_1320_n66# a_1106_n54302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14960 word409 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14961 GND A0 word1012 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14962 word635 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14963 a_2162_n98748# a_2112_n66# a_1898_n98748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14964 word883 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14965 a_1898_n136378# a_1848_n66# a_1634_n136378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14966 word748 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14967 a_578_n100026# a_528_n66# a_446_n100026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14968 a_1370_n103434# a_1320_n66# a_1238_n103434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14969 a_1898_n128000# a_1848_n66# a_1766_n128000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14970 a_446_n19228# A8 a_182_n19228# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14971 GND A7 word111 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14972 a_1766_n23772# A3 a_1502_n23772# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14973 GND A7 word60 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14974 word569 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14975 word981 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14976 GND A5 word712 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14977 word538 A0 a_2162_n76596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14978 GND A7 word885 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14979 GND A9 word26 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14980 a_578_n138508# a_528_n66# a_314_n138508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14981 GND A9 word354 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14982 word947 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14983 word44 A0 a_2294_n6448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14984 a_446_n88524# A8 a_50_n88524# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14985 a_2294_n126864# A1 a_1898_n126864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14986 GND A5 word200 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14987 a_1106_n9146# a_1056_n66# a_974_n9146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14988 word93 a_2376_n66# a_2294_n13406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14989 word104 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X14990 a_2294_n96760# A1 a_2030_n96760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14991 word877 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14992 word936 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14993 GND A1 word1008 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14994 GND A1 word949 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14995 word675 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14996 word953 a_2376_n66# a_2294_n135526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X14997 GND A4 word806 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14998 a_446_n10140# A8 a_182_n10140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X14999 a_2030_n84264# A2 a_1766_n84264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15000 GND A8 word524 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15001 word917 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15002 a_1370_n22352# a_1320_n66# a_1238_n22352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15003 word651 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15004 word725 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15005 word1002 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15006 word955 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15007 GND A0 word846 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15008 a_1766_n39108# A3 a_1370_n39108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15009 GND A8 word92 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15010 GND A7 word377 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15011 word581 a_2376_n66# a_2294_n82702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15012 a_1766_n61544# A3 a_1370_n61544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15013 a_446_n106274# A8 a_50_n106274# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15014 GND A1 word517 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15015 a_1238_n109682# A5 a_974_n109682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15016 word65 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15017 a_710_n79294# A7 a_446_n79294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15018 GND A6 word21 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15019 a_1238_n101020# A5 a_842_n101020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15020 word756 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15021 a_1106_n42516# a_1056_n66# a_974_n42516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15022 a_578_n106558# a_528_n66# a_446_n106558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15023 a_2030_n113090# A2 a_1634_n113090# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15024 word429 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15025 a_710_n115220# A7 a_314_n115220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15026 GND A2 word641 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15027 GND A9 word459 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15028 a_1502_n118628# A4 a_1238_n118628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15029 a_2294_n1904# A1 a_1898_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15030 a_1766_n30020# A3 a_1370_n30020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15031 GND A9 word400 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15032 a_1238_n100594# A5 a_842_n100594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15033 word268 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15034 word139 a_2376_n66# a_2162_n19938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15035 word426 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15036 word982 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15037 a_446_n25050# A8 a_182_n25050# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15038 a_2030_n99174# A2 a_1634_n99174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15039 word730 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15040 GND A4 word911 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15041 GND A1 word20 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15042 a_710_n114794# A7 a_314_n114794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15043 a_1370_n98606# a_1320_n66# a_1106_n98606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15044 a_710_n123172# A7 a_314_n123172# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15045 GND A1 word292 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15046 word1022 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15047 GND A8 word629 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15048 GND A2 word360 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15049 a_1106_n71910# a_1056_n66# a_842_n71910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15050 GND A7 word541 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15051 GND A0 word892 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15052 a_578_n144330# a_528_n66# a_314_n144330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15053 GND A8 word138 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15054 GND A8 word197 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15055 word60 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15056 a_446_n85968# A8 a_50_n85968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15057 a_446_n94346# A8 a_50_n94346# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15058 a_2294_n141064# A1 a_2030_n141064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15059 a_2294_n132686# A1 a_1898_n132686# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15060 a_974_n41806# A6 a_710_n41806# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15061 word918 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15062 GND A3 word994 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15063 a_1106_n6590# a_1056_n66# a_974_n6590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15064 word75 a_2376_n66# a_2162_n10850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15065 GND A3 word935 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15066 GND A4 word847 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15067 a_2030_n90086# A2 a_1634_n90086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15068 word935 a_2376_n66# a_2162_n132970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15069 a_710_n4744# A7 a_446_n4744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15070 word475 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15071 GND A8 word565 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15072 word405 a_2376_n66# a_2294_n57710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15073 GND A7 word260 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15074 a_842_n11844# a_792_n66# a_710_n11844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15075 a_974_n18944# A6 a_578_n18944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15076 a_974_n27322# A6 a_578_n27322# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15077 word816 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15078 GND A1 word888 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15079 GND A3 word833 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15080 word833 a_2376_n66# a_2294_n118486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15081 a_1370_n66656# a_1320_n66# a_1238_n66656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15082 word797 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15083 GND A0 word726 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15084 word894 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15085 a_1898_n5312# a_1848_n66# a_1766_n5312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15086 word461 a_2376_n66# a_2294_n65662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15087 GND A7 word316 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15088 a_50_n114652# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15089 word312 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15090 GND A1 word397 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15091 GND A7 word257 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15092 a_1106_n86820# a_1056_n66# a_842_n86820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15093 GND A5 word858 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15094 GND A2 word465 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15095 GND A9 word500 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15096 a_1502_n124450# A4 a_1106_n124450# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15097 GND A5 word799 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15098 a_1106_n25476# a_1056_n66# a_974_n25476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15099 GND A6 word156 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15100 word250 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15101 a_974_n56716# A6 a_578_n56716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15102 word239 a_2376_n66# a_2162_n34138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15103 word1023 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15104 GND A0 word158 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15105 GND A2 word521 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15106 word829 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15107 GND A8 word670 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15108 a_842_n35132# a_792_n66# a_578_n35132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15109 GND A0 word992 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15110 word51 a_2376_n66# a_2162_n7442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15111 GND A7 word523 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15112 GND A8 word740 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15113 word781 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15114 a_446_n91790# A8 a_50_n91790# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15115 a_1766_n82276# A3 a_1502_n82276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15116 GND A1 word604 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15117 GND A0 word646 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15118 a_182_n16104# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15119 word87 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15120 GND A4 word481 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15121 a_1766_n73898# A3 a_1502_n73898# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15122 GND A2 word240 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15123 a_1106_n63248# a_1056_n66# a_974_n63248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15124 GND A6 word422 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15125 a_1370_n139076# a_1320_n66# a_1238_n139076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15126 word767 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15127 a_1370_n4602# a_1320_n66# a_1238_n4602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15128 a_1898_n37404# a_1848_n66# a_1766_n37404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15129 a_446_n6164# A8 a_182_n6164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15130 a_50_n129562# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15131 GND A5 word904 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15132 GND A6 word693 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15133 a_974_n24766# A6 a_578_n24766# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15134 word141 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15135 GND A6 word261 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15136 GND A0 word424 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15137 GND A2 word986 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15138 a_2162_n2188# a_2112_n66# a_1898_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15139 word636 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15140 word62 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15141 a_50_n85542# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15142 a_842_n64526# a_792_n66# a_578_n64526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15143 word412 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15144 a_1370_n72478# a_1320_n66# a_1106_n72478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15145 a_2294_n8152# A1 a_2030_n8152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15146 word143 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15147 GND A2 word626 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15148 word703 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15149 a_50_n120474# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15150 a_1502_n27606# A4 a_1238_n27606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15151 GND A4 word256 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15152 GND A2 word705 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15153 word287 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15154 word974 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15155 word886 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15156 word624 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15157 GND A7 word628 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15158 a_578_n23346# a_528_n66# a_446_n23346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15159 a_842_n103434# a_792_n66# a_578_n103434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15160 a_1502_n96902# A4 a_1106_n96902# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15161 GND A3 word96 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15162 a_974_n62538# A6 a_578_n62538# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15163 a_1106_n78158# a_1056_n66# a_974_n78158# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15164 GND A2 word345 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15165 a_1106_n69780# a_1056_n66# a_842_n69780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15166 GND A6 word527 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15167 a_578_n92642# a_528_n66# a_446_n92642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15168 word929 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15169 word870 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15170 a_314_n43510# a_264_n66# a_182_n43510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15171 GND A4 word39 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15172 word246 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15173 word119 a_2376_n66# a_2162_n17098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15174 a_842_n32576# a_792_n66# a_578_n32576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15175 a_974_n39676# A6 a_710_n39676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15176 GND A0 word470 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15177 GND A7 word564 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15178 a_1766_n3466# A3 a_1370_n3466# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15179 word33 a_2376_n66# a_2294_n4886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15180 GND A1 word645 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15181 GND A4 word463 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15182 GND A4 word522 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15183 a_182_n13548# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15184 a_314_n51462# a_264_n66# a_182_n51462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15185 word248 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15186 GND A8 word550 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15187 word86 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15188 a_578_n61118# a_528_n66# a_314_n61118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15189 a_1898_n43226# a_1848_n66# a_1634_n43226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15190 a_842_n141206# a_792_n66# a_578_n141206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15191 a_842_n18092# a_792_n66# a_710_n18092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15192 a_1898_n34848# a_1848_n66# a_1766_n34848# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15193 word607 a_2376_n66# a_2162_n86394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15194 a_50_n135384# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15195 GND A0 word526 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15196 a_1502_n64952# A4 a_1238_n64952# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15197 a_314_n144614# a_264_n66# a_50_n144614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15198 word451 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15199 word392 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15200 GND A2 word810 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15201 a_1634_n20506# a_1584_n66# a_1502_n20506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15202 GND A6 word302 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15203 a_842_n118344# a_792_n66# a_710_n118344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15204 a_578_n29878# a_528_n66# a_446_n29878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15205 word44 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15206 a_578_n60692# a_528_n66# a_314_n60692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15207 a_182_n59982# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15208 a_50_n82986# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15209 a_50_n91364# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15210 a_842_n70348# a_792_n66# a_578_n70348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15211 word453 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15212 a_974_n77448# A6 a_710_n77448# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15213 a_1634_n4176# a_1584_n66# a_1370_n4176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15214 GND A0 word304 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15215 GND A2 word866 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15216 a_182_n51320# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15217 a_314_n58420# a_264_n66# a_182_n58420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15218 GND A2 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15219 a_1502_n33428# A4 a_1106_n33428# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15220 word516 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15221 GND A4 word297 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15222 word455 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15223 GND A4 word238 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15224 a_1898_n72620# a_1848_n66# a_1634_n72620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15225 word1015 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15226 a_1238_n2756# A5 a_974_n2756# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15227 a_842_n47486# a_792_n66# a_710_n47486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15228 word665 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15229 word960 A0 a_2294_n136520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15230 word868 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15231 a_1766_n9998# A3 a_1502_n9998# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15232 a_1898_n11276# a_1848_n66# a_1634_n11276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15233 a_842_n100878# a_792_n66# a_578_n100878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15234 a_182_n28458# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15235 a_578_n20790# a_528_n66# a_446_n20790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15236 a_1238_n10708# A5 a_842_n10708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15237 a_314_n57994# a_264_n66# a_182_n57994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15238 a_314_n66372# a_264_n66# a_182_n66372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15239 a_314_n121042# a_264_n66# a_50_n121042# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15240 a_182_n50894# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15241 word191 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15242 a_314_n112664# a_264_n66# a_50_n112664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15243 word511 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15244 a_578_n67650# a_528_n66# a_314_n67650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15245 a_1898_n49758# a_1848_n66# a_1634_n49758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15246 a_1502_n1052# A4 a_1238_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15247 a_2030_n8294# A2 a_1634_n8294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15248 GND A3 word49 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15249 word59 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15250 GND A3 word467 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15251 a_1898_n80572# a_1848_n66# a_1766_n80572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15252 word1016 A0 a_2294_n144472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15253 word660 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15254 a_1766_n125302# A3 a_1370_n125302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15255 a_1766_n116924# A3 a_1370_n116924# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15256 word193 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15257 GND A0 word570 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15258 a_974_n113516# A6 a_710_n113516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15259 word228 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15260 a_1634_n35416# a_1584_n66# a_1370_n35416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15261 a_974_n45498# A6 a_710_n45498# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15262 word1001 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15263 word942 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15264 word809 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15265 a_182_n1194# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15266 word39 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15267 word750 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15268 a_2162_n111812# a_2112_n66# a_2030_n111812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15269 a_50_n97896# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15270 a_842_n85258# a_792_n66# a_710_n85258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15271 word558 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15272 a_2162_n26612# a_2112_n66# a_2030_n26612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15273 word230 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15274 word790 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15275 a_182_n66230# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15276 word126 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15277 a_1898_n40670# a_1848_n66# a_1634_n40670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15278 GND A0 word350 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15279 word499 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15280 GND A2 word971 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15281 word462 A0 a_2162_n65804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15282 word440 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15283 word621 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15284 word398 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15285 word492 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15286 word275 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15287 a_1898_n87530# a_1848_n66# a_1766_n87530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15288 word720 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15289 word433 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15290 word128 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15291 word973 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15292 a_842_n124166# a_792_n66# a_710_n124166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15293 a_578_n35700# a_528_n66# a_446_n35700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15294 a_1898_n26186# a_1848_n66# a_1766_n26186# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15295 GND A3 word674 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15296 word338 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15297 GND A3 word242 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15298 word494 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15299 GND A9 word117 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15300 a_2294_n24624# A1 a_1898_n24624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15301 a_314_n127574# a_264_n66# a_50_n127574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15302 a_1898_n95482# a_1848_n66# a_1634_n95482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15303 a_1238_n94914# A5 a_974_n94914# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15304 word776 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15305 a_1898_n102014# a_1848_n66# a_1634_n102014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15306 a_974_n128426# A6 a_578_n128426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15307 word333 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15308 word110 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15309 word456 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15310 a_1634_n72762# a_1584_n66# a_1370_n72762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15311 a_2162_n126722# a_2112_n66# a_2030_n126722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15312 a_182_n34280# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15313 word296 A0 a_2294_n42232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15314 GND A4 word609 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15315 a_314_n72194# a_264_n66# a_182_n72194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15316 word394 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15317 a_1634_n122462# a_1584_n66# a_1370_n122462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15318 word895 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15319 a_1898_n55580# a_1848_n66# a_1766_n55580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15320 word840 A0 a_2294_n119480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15321 word166 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15322 GND A3 word449 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15323 GND A6 word787 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15324 word234 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15325 a_974_n110960# A6 a_710_n110960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15326 word825 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15327 a_2030_n41522# A2 a_1766_n41522# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15328 word315 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15329 a_842_n139076# a_792_n66# a_578_n139076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15330 a_1370_n8294# a_1320_n66# a_1106_n8294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15331 word848 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15332 a_1898_n131408# a_1848_n66# a_1634_n131408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15333 a_2294_n39534# A1 a_1898_n39534# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15334 word540 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15335 word599 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15336 a_974_n98180# A6 a_578_n98180# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15337 a_2162_n32434# a_2112_n66# a_2030_n32434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15338 a_710_n36552# A7 a_314_n36552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15339 GND A0 word450 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15340 word562 A0 a_2162_n80004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15341 word371 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15342 a_1634_n129420# a_1584_n66# a_1502_n129420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15343 word746 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15344 word439 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15345 word169 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15346 word701 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15347 word1014 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15348 a_446_n13832# A8 a_182_n13832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15349 a_1238_n31440# A5 a_842_n31440# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15350 word432 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15351 a_1634_n87672# a_1584_n66# a_1502_n87672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15352 a_182_n49190# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15353 word342 A0 a_2162_n48764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15354 GND A9 word217 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15355 GND A9 word158 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15356 a_2030_n117208# A2 a_1634_n117208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15357 a_314_n133396# a_264_n66# a_50_n133396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15358 word751 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15359 a_1106_n145182# a_1056_n66# a_842_n145182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15360 a_2294_n30446# A1 a_1898_n30446# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15361 word278 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15362 a_2030_n70916# A2 a_1766_n70916# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15363 word657 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15364 a_1634_n128994# a_1584_n66# a_1502_n128994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15365 word149 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15366 GND A5 word653 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15367 GND A5 word221 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15368 GND A3 word613 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15369 GND A6 word951 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15370 a_2162_n61828# a_2112_n66# a_2030_n61828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15371 a_2294_n68928# A1 a_1898_n68928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15372 word339 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15373 a_446_n101304# A8 a_50_n101304# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15374 a_974_n134248# A6 a_578_n134248# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15375 GND A1 word812 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15376 a_1634_n56148# a_1584_n66# a_1502_n56148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15377 a_710_n74324# A7 a_446_n74324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15378 word479 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15379 a_1634_n47770# a_1584_n66# a_1502_n47770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15380 word497 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15381 word120 A0 a_2294_n17240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15382 a_1238_n86252# A5 a_842_n86252# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15383 word637 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15384 GND A4 word650 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15385 a_1106_n105280# a_1056_n66# a_842_n105280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15386 a_710_n118912# A7 a_314_n118912# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15387 word214 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15388 a_1502_n69070# A4 a_1106_n69070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15389 word639 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15390 word608 A0 a_2294_n86536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15391 GND A9 word424 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15392 word1017 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15393 word176 A0 a_2294_n25192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15394 a_2162_n109682# a_2112_n66# a_2030_n109682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15395 a_2030_n16530# A2 a_1766_n16530# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15396 GND A5 word270 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15397 a_2162_n101020# a_2112_n66# a_1898_n101020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15398 a_446_n28742# A8 a_182_n28742# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15399 word174 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15400 a_1238_n46350# A5 a_842_n46350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15401 word605 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15402 GND A3 word388 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15403 GND A9 word263 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15404 a_1766_n114084# A3 a_1502_n114084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15405 word114 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15406 a_2030_n85826# A2 a_1634_n85826# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15407 a_710_n42374# A7 a_314_n42374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15408 a_1634_n24198# a_1584_n66# a_1502_n24198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15409 a_2030_n24482# A2 a_1634_n24482# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15410 word195 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15411 GND A5 word326 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15412 GND A8 word162 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15413 a_2162_n85116# a_2112_n66# a_1898_n85116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15414 GND A8 word103 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15415 a_2162_n76738# a_2112_n66# a_2030_n76738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15416 a_2162_n100594# a_2112_n66# a_2030_n100594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15417 word728 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15418 a_1238_n119622# A5 a_842_n119622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15419 a_1898_n114368# a_1848_n66# a_1766_n114368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15420 a_710_n89234# A7 a_446_n89234# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15421 a_446_n107836# A8 a_50_n107836# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15422 word602 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15423 a_2162_n15394# a_2112_n66# a_2030_n15394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15424 GND A1 word96 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15425 GND A6 word32 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15426 GND A7 word789 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15427 word911 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15428 a_2030_n123030# A2 a_1766_n123030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15429 a_1634_n143194# a_1584_n66# a_1502_n143194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15430 word851 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15431 word319 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15432 a_1766_n48622# A3 a_1370_n48622# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15433 a_2294_n113232# A1 a_1898_n113232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15434 word51 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15435 a_2294_n104854# A1 a_2030_n104854# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15436 GND A3 word595 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15437 GND A6 word933 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15438 GND A9 word470 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15439 word380 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15440 a_2294_n74750# A1 a_1898_n74750# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15441 a_2294_n83128# A1 a_2030_n83128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15442 a_1238_n110534# A5 a_974_n110534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15443 word781 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15444 a_1766_n143478# A3 a_1370_n143478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15445 GND A1 word853 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15446 a_710_n80146# A7 a_446_n80146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15447 a_2030_n53876# A2 a_1634_n53876# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15448 GND A5 word592 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15449 GND A5 word533 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15450 a_1238_n92074# A5 a_974_n92074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15451 word994 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15452 a_1238_n83696# A5 a_842_n83696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15453 a_710_n910# A7 a_446_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15454 GND A2 word491 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15455 GND A7 word281 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15456 a_710_n124734# A7 a_314_n124734# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15457 a_2162_n44788# a_2112_n66# a_2030_n44788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15458 GND A8 word47 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15459 a_1370_n38824# a_1320_n66# a_1238_n38824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15460 GND A8 word208 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15461 word590 A0 a_2162_n83980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15462 word833 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15463 GND A0 word962 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15464 a_1898_n129278# a_1848_n66# a_1634_n129278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15465 a_446_n95908# A8 a_50_n95908# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15466 word856 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15467 GND A1 word201 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15468 a_446_n34564# A8 a_182_n34564# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15469 a_1766_n16672# A3 a_1370_n16672# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15470 GND A7 word835 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15471 GND A7 word894 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15472 word488 A0 a_2294_n69496# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15473 GND A9 word304 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15474 GND A2 word427 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15475 GND A9 word245 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15476 word1005 a_2376_n66# a_2294_n142910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15477 word897 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15478 a_2294_n42800# A1 a_1898_n42800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15479 GND A8 word766 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15480 a_2294_n128142# A1 a_1898_n128142# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15481 word295 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15482 a_2294_n98038# A1 a_2030_n98038# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15483 GND A8 word705 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15484 word886 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15485 a_2162_n6306# a_2112_n66# a_2030_n6306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15486 GND A7 word66 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15487 GND A8 word144 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15488 word485 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15489 word827 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15490 GND A3 word903 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15491 a_1898_n120190# a_1848_n66# a_1634_n120190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15492 GND A2 word266 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15493 word903 a_2376_n66# a_2162_n128426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15494 a_2030_n68786# A2 a_1766_n68786# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15495 a_710_n86678# A7 a_446_n86678# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15496 word601 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15497 a_2162_n144898# a_2112_n66# a_2030_n144898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15498 word531 a_2376_n66# a_2162_n75602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15499 word952 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15500 word905 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15501 a_1370_n125728# a_1320_n66# a_1106_n125728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15502 GND A0 word796 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15503 a_2162_n59698# a_2112_n66# a_2030_n59698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15504 a_2162_n68076# a_2112_n66# a_1898_n68076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15505 GND A7 word327 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15506 a_974_n8436# A6 a_710_n8436# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15507 word33 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15508 a_1106_n35416# a_1056_n66# a_842_n35416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15509 GND A6 word167 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15510 word690 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15511 a_578_n130272# a_528_n66# a_314_n130272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15512 word379 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15513 word683 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15514 GND A7 word105 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15515 GND A9 word409 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15516 GND A9 word350 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15517 a_2294_n66088# A1 a_2030_n66088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15518 GND A1 word733 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15519 a_1502_n142342# A4 a_1106_n142342# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15520 GND A4 word963 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15521 a_1502_n133964# A4 a_1106_n133964# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15522 GND A9 word20 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15523 a_1370_n53024# a_1320_n66# a_1106_n53024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15524 a_1370_n44646# a_1320_n66# a_1106_n44646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15525 GND A8 word249 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15526 GND A7 word593 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15527 word376 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15528 a_1898_n135100# a_1848_n66# a_1766_n135100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15529 a_710_n116072# A7 a_314_n116072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15530 GND A7 word102 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15531 word913 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15532 GND A0 word842 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15533 a_578_n137230# a_528_n66# a_314_n137230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15534 a_50_n139502# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15535 a_446_n87246# A8 a_50_n87246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15536 a_446_n7726# A8 a_182_n7726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15537 a_446_n78868# A8 a_50_n78868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15538 a_1766_n69354# A3 a_1502_n69354# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15539 GND A5 word974 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15540 word95 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15541 word154 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15542 GND A6 word272 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15543 word868 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15544 GND A3 word944 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15545 GND A1 word940 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15546 a_1238_n131266# A5 a_974_n131266# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15547 GND A3 word885 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15548 GND A2 word307 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15549 a_1106_n72762# a_1056_n66# a_842_n72762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15550 word885 a_2376_n66# a_2294_n125870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15551 a_578_n145182# a_528_n66# a_314_n145182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15552 a_1502_n110392# A4 a_1238_n110392# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15553 a_710_n6022# A7 a_446_n6022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15554 GND A4 word738 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15555 GND A8 word515 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15556 word849 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15557 a_842_n13122# a_792_n66# a_710_n13122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15558 a_1370_n12696# a_1320_n66# a_1238_n12696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15559 a_1370_n21074# a_1320_n66# a_1238_n21074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15560 GND A2 word696 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15561 a_1370_n131550# a_1320_n66# a_1238_n131550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15562 GND A0 word778 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15563 a_50_n130414# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15564 GND A7 word368 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15565 a_1766_n60266# A3 a_1502_n60266# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15566 GND A1 word449 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15567 GND A1 word508 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15568 a_974_n5880# A6 a_710_n5880# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15569 a_1106_n41238# a_1056_n66# a_974_n41238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15570 a_1106_n32860# a_1056_n66# a_842_n32860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15571 word411 a_2376_n66# a_2162_n58562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15572 a_578_n105280# a_528_n66# a_446_n105280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15573 a_1766_n98748# A3 a_1370_n98748# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15574 a_1370_n108688# a_1320_n66# a_1106_n108688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15575 GND A8 word571 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15576 a_1370_n117066# a_1320_n66# a_1106_n117066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15577 a_578_n24908# a_528_n66# a_446_n24908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15578 word1002 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15579 a_50_n107552# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15580 a_1106_n79720# a_1056_n66# a_974_n79720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15581 GND A9 word450 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15582 GND A4 word1004 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15583 word719 a_2376_n66# a_2162_n102298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15584 word189 a_2376_n66# a_2294_n27038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15585 word200 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15586 GND A7 word634 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15587 a_1106_n87672# a_1056_n66# a_842_n87672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15588 GND A7 word575 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15589 word914 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15590 word973 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15591 a_1238_n137798# A5 a_842_n137798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15592 a_182_n5312# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15593 GND A0 word108 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15594 GND A4 word902 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15595 a_314_n61402# a_264_n66# a_182_n61402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15596 a_1370_n88950# a_1320_n66# a_1106_n88950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15597 word1013 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15598 word996 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15599 GND A8 word620 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15600 GND A4 word101 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15601 word954 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15602 a_842_n28032# a_792_n66# a_578_n28032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15603 word677 a_2376_n66# a_2294_n96334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15604 a_50_n136946# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15605 a_50_n145324# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15606 a_446_n93068# A8 a_50_n93068# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15607 GND A0 word596 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15608 GND A1 word613 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15609 a_446_n84690# A8 a_50_n84690# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15610 a_1766_n66798# A3 a_1370_n66798# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15611 a_1766_n75176# A3 a_1370_n75176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15612 word462 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15613 a_974_n40528# A6 a_710_n40528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15614 GND A6 word313 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15615 GND A8 word676 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15616 a_842_n119906# a_792_n66# a_710_n119906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15617 a_578_n70632# a_528_n66# a_314_n70632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15618 word850 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15619 word985 a_2376_n66# a_2294_n140070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15620 a_710_n3466# A7 a_446_n3466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15621 a_182_n69922# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15622 a_50_n92926# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15623 a_842_n71910# a_792_n66# a_578_n71910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15624 a_974_n26044# A6 a_578_n26044# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15625 GND A0 word374 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15626 GND A2 word936 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15627 a_842_n10566# a_792_n66# a_710_n10566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15628 GND A4 word367 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15629 word586 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15630 a_50_n78442# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15631 a_1370_n57000# a_1320_n66# a_1238_n57000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15632 word788 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15633 a_1898_n21216# a_1848_n66# a_1766_n21216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15634 a_578_n30730# a_528_n66# a_446_n30730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15635 a_50_n113374# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15636 a_50_n104996# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15637 word244 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15638 GND A1 word388 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15639 a_182_n60834# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15640 a_314_n67934# a_264_n66# a_182_n67934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15641 GND A4 word206 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15642 a_1502_n42942# A4 a_1106_n42942# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15643 a_314_n122604# a_264_n66# a_50_n122604# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15644 word296 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15645 GND A5 word790 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15646 a_1106_n24198# a_1056_n66# a_974_n24198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15647 GND A6 word147 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15648 a_1898_n90512# a_1848_n66# a_1634_n90512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15649 a_446_n99600# A8 a_50_n99600# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15650 a_182_n37972# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15651 a_974_n55438# A6 a_578_n55438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15652 GND A6 word418 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15653 word1014 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15654 word1012 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15655 word879 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15656 GND A0 word90 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15657 word820 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15658 a_182_n2756# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15659 a_1502_n11418# A4 a_1238_n11418# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15660 a_710_n9998# A7 a_446_n9998# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15661 GND A4 word142 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15662 a_842_n86820# a_792_n66# a_710_n86820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15663 word196 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15664 GND A0 word420 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15665 word659 a_2376_n66# a_2162_n93778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15666 GND A7 word514 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15667 a_50_n142768# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15668 word510 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15669 word691 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15670 word632 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15671 word503 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15672 word876 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15673 a_314_n44362# a_264_n66# a_182_n44362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15674 word139 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15675 word198 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15676 a_446_n200# A8 a_182_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15677 a_1370_n3324# a_1320_n66# a_1238_n3324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15678 a_1502_n10992# A4 a_1238_n10992# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15679 a_1898_n36126# a_1848_n66# a_1634_n36126# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15680 word557 a_2376_n66# a_2294_n79294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15681 a_842_n125728# a_792_n66# a_710_n125728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15682 a_50_n128284# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15683 word349 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15684 word408 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15685 GND A0 word476 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15686 a_974_n93210# A6 a_578_n93210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15687 word566 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15688 a_314_n137514# a_264_n66# a_50_n137514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15689 GND A6 word684 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15690 word686 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15691 word401 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15692 GND A2 word760 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15693 word342 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15694 a_1634_n13406# a_1584_n66# a_1370_n13406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15695 a_974_n23488# A6 a_578_n23488# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15696 word846 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15697 word787 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15698 word568 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15699 a_50_n84264# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15700 a_1370_n71200# a_1320_n66# a_1106_n71200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15701 a_50_n75886# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15702 a_974_n92784# A6 a_578_n92784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15703 GND A2 word816 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15704 a_182_n44220# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15705 GND A0 word254 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15706 GND A4 word679 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15707 GND A2 word43 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15708 word285 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15709 word243 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15710 word405 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15711 a_1238_n4034# A5 a_974_n4034# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15712 a_1898_n65520# a_1848_n66# a_1634_n65520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15713 GND A7 word619 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15714 a_842_n102156# a_792_n66# a_578_n102156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15715 GND A1 word700 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15716 word910 A0 a_2162_n129420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15717 word759 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15718 a_578_n22068# a_528_n66# a_446_n22068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15719 word183 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15720 word236 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15721 a_1502_n95624# A4 a_1106_n95624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15722 a_314_n59272# a_264_n66# a_182_n59272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15723 a_182_n43794# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15724 a_182_n52172# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15725 GND A3 word87 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15726 a_974_n61260# A6 a_578_n61260# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15727 a_1106_n108972# a_1056_n66# a_842_n108972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15728 a_2030_n111812# A2 a_1766_n111812# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15729 GND A6 word400 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15730 word461 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15731 GND A3 word417 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15732 a_1898_n73472# a_1848_n66# a_1766_n73472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15733 a_578_n91364# a_528_n66# a_446_n91364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15734 a_1238_n72904# A5 a_974_n72904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15735 word671 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15736 word966 A0 a_2162_n137372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15737 a_1766_n109824# A3 a_1502_n109824# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15738 a_974_n38398# A6 a_710_n38398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15739 GND A0 word520 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15740 a_1634_n19938# a_1584_n66# a_1502_n19938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15741 a_842_n31298# a_792_n66# a_578_n31298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15742 word441 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15743 word951 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15744 word892 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15745 GND A4 word513 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15746 word673 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15747 a_182_n12270# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15748 a_50_n99174# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15749 GND A0 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15750 GND A4 word454 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15751 a_314_n50184# a_264_n66# a_182_n50184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15752 word82 A0 a_2162_n11844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15753 a_842_n69780# a_792_n66# a_578_n69780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15754 word180 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15755 word239 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15756 word631 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15757 a_1898_n140922# a_1848_n66# a_1634_n140922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15758 a_1634_n97612# a_1584_n66# a_1502_n97612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15759 a_182_n59130# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15760 word412 A0 a_2294_n58704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15761 GND A3 word294 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15762 GND A3 word353 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15763 word79 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15764 a_314_n134958# a_264_n66# a_50_n134958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15765 a_314_n143336# a_264_n66# a_50_n143336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15766 a_1766_n100736# A3 a_1502_n100736# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15767 word383 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15768 a_1634_n10850# a_1584_n66# a_1502_n10850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15769 a_1898_n19086# a_1848_n66# a_1766_n19086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15770 GND A3 word624 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15771 a_578_n28600# a_528_n66# a_446_n28600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15772 a_1238_n18518# A5 a_974_n18518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15773 a_842_n108688# a_792_n66# a_578_n108688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15774 a_182_n67082# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15775 a_50_n90086# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15776 GND A3 word192 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15777 a_1238_n40954# A5 a_974_n40954# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15778 a_974_n135810# A6 a_578_n135810# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15779 a_974_n76170# A6 a_710_n76170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15780 word444 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15781 a_2030_n126722# A2 a_1634_n126722# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15782 a_710_n14542# A7 a_446_n14542# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15783 word76 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15784 a_578_n97896# a_528_n66# a_446_n97896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15785 a_1898_n88382# a_1848_n66# a_1634_n88382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15786 word726 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15787 a_1106_n115220# a_1056_n66# a_974_n115220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15788 GND A2 word25 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15789 a_1502_n32150# A4 a_1106_n32150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15790 GND A4 word288 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15791 a_2162_n48906# a_2112_n66# a_1898_n48906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15792 a_1502_n79010# A4 a_1106_n79010# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15793 a_1238_n1478# A5 a_974_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15794 a_1634_n65662# a_1584_n66# a_1502_n65662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15795 GND A4 word559 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15796 a_182_n27180# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15797 a_314_n65094# a_264_n66# a_182_n65094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15798 word246 A0 a_2162_n35132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15799 word182 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15800 a_314_n111386# a_264_n66# a_50_n111386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15801 a_1106_n123172# a_1056_n66# a_842_n123172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15802 a_1634_n115362# a_1584_n66# a_1502_n115362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15803 a_1106_n114794# a_1056_n66# a_974_n114794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15804 word123 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15805 a_1898_n48480# a_1848_n66# a_1766_n48480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15806 word502 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15807 word50 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15808 word116 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15809 a_1502_n78584# A4 a_1106_n78584# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15810 GND A6 word796 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15811 a_2294_n46918# A1 a_2030_n46918# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15812 a_974_n112238# A6 a_710_n112238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15813 word488 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15814 a_1634_n34138# a_1584_n66# a_1502_n34138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15815 word125 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15816 a_710_n52314# A7 a_314_n52314# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15817 GND A8 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15818 word611 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15819 word992 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15820 a_710_n43936# A7 a_314_n43936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15821 a_2030_n34422# A2 a_1766_n34422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15822 word265 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15823 GND A5 word396 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15824 word933 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15825 word30 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15826 a_1238_n64242# A5 a_842_n64242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15827 a_1238_n55864# A5 a_974_n55864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15828 GND A4 word495 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15829 word549 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15830 a_1898_n115930# a_1848_n66# a_1634_n115930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15831 a_1766_n11702# A3 a_1370_n11702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15832 a_2162_n16956# a_2112_n66# a_1898_n16956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15833 a_1502_n47060# A4 a_1238_n47060# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15834 word981 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15835 word321 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15836 a_314_n140780# a_264_n66# a_50_n140780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15837 a_1634_n144756# a_1584_n66# a_1370_n144756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15838 word964 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15839 a_1898_n123882# a_1848_n66# a_1766_n123882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15840 word382 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15841 GND A2 a_1848_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X15842 GND A7 word31 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15843 GND A7 word856 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15844 GND A9 word108 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15845 a_710_n81708# A7 a_446_n81708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15846 a_2030_n63816# A2 a_1766_n63816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15847 a_314_n126296# a_264_n66# a_50_n126296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15848 GND A5 word662 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15849 a_2294_n14968# A1 a_2030_n14968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15850 GND A5 word603 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15851 word99 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15852 a_1238_n93636# A5 a_974_n93636# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15853 GND A6 word901 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15854 word1005 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15855 word917 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15856 a_710_n11986# A7 a_446_n11986# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15857 a_2162_n63106# a_2112_n66# a_2030_n63106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15858 a_1634_n49048# a_1584_n66# a_1370_n49048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15859 a_2030_n49332# A2 a_1634_n49332# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15860 word506 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15861 a_2030_n109682# A2 a_1766_n109682# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15862 word587 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15863 word660 A0 a_2294_n93920# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15864 word655 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15865 a_2162_n125444# a_2112_n66# a_2030_n125444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15866 word228 A0 a_2294_n32576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15867 word756 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15868 GND A3 word499 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15869 word558 A0 a_2162_n79436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15870 GND A9 word374 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15871 GND A9 word46 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15872 a_2294_n61118# A1 a_1898_n61118# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15873 GND A9 word315 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15874 word967 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15875 GND A6 word778 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15876 word126 A0 a_2162_n18092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15877 word225 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15878 a_1766_n121468# A3 a_1370_n121468# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15879 word365 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15880 a_2030_n100594# A2 a_1766_n100594# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15881 a_2294_n129704# A1 a_2030_n129704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15882 word124 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15883 a_2030_n40244# A2 a_1634_n40244# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15884 word487 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15885 a_1238_n39250# A5 a_974_n39250# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15886 GND A3 word338 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15887 a_2294_n29878# A1 a_2030_n29878# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15888 a_2162_n31156# a_2112_n66# a_2030_n31156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15889 a_2294_n38256# A1 a_1898_n38256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15890 GND A2 word336 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15891 a_2030_n78726# A2 a_1634_n78726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15892 a_710_n111102# A7 a_314_n111102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15893 GND A9 word371 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15894 a_2162_n22778# a_2112_n66# a_1898_n22778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15895 a_1370_n16814# a_1320_n66# a_1106_n16814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15896 a_2030_n17382# A2 a_1634_n17382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15897 word494 A0 a_2162_n70348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15898 word1022 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15899 GND A5 word276 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15900 GND A8 word112 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15901 word963 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15902 word430 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15903 a_446_n109114# A8 a_50_n109114# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15904 a_2294_n120616# A1 a_2030_n120616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15905 a_446_n12554# A8 a_182_n12554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15906 GND A6 word41 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15907 word423 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15908 a_1634_n86394# a_1584_n66# a_1370_n86394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15909 word364 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15910 GND A9 word149 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15911 GND A9 word90 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15912 a_1634_n136094# a_1584_n66# a_1370_n136094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15913 a_578_n140212# a_528_n66# a_314_n140212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15914 a_578_n131834# a_528_n66# a_314_n131834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15915 a_5140_164# A8 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X15916 a_2294_n20790# A1 a_2030_n20790# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15917 GND A5 word644 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15918 word694 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15919 word31 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15920 GND A9 word479 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15921 GND A3 word545 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15922 GND A9 word420 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15923 word330 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15924 a_446_n100026# A8 a_50_n100026# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15925 a_1238_n103434# A5 a_842_n103434# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15926 GND A1 word744 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15927 a_1766_n128000# A3 a_1502_n128000# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15928 a_2030_n55154# A2 a_1766_n55154# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15929 a_710_n73046# A7 a_446_n73046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15930 a_2030_n46776# A2 a_1634_n46776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15931 a_578_n108972# a_528_n66# a_446_n108972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15932 GND A5 word542 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15933 word446 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15934 word569 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15935 word885 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15936 a_1898_n145040# a_1848_n66# a_1634_n145040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15937 a_2162_n131266# a_2112_n66# a_2030_n131266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15938 a_1238_n76596# A5 a_974_n76596# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15939 a_578_n100310# a_528_n66# a_446_n100310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15940 a_1370_n103718# a_1320_n66# a_1238_n103718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15941 word738 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15942 a_710_n126012# A7 a_314_n126012# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15943 a_2162_n46066# a_2112_n66# a_2030_n46066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15944 a_710_n117634# A7 a_314_n117634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15945 GND A9 word476 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15946 a_1766_n32434# A3 a_1502_n32434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15947 GND A1 word312 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15948 GND A8 word56 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15949 GND A0 word912 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15950 word540 A0 a_2294_n76880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15951 a_446_n88808# A8 a_50_n88808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15952 word535 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15953 a_2294_n135526# A1 a_2030_n135526# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15954 word949 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15955 a_446_n27464# A8 a_182_n27464# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15956 GND A1 word37 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15957 GND A2 word377 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15958 GND A9 word254 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15959 GND A9 word195 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15960 GND A4 word867 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15961 a_2294_n44078# A1 a_1898_n44078# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15962 a_2030_n84548# A2 a_1766_n84548# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15963 a_2030_n144898# A2 a_1634_n144898# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15964 word955 a_2376_n66# a_2162_n135810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15965 a_1502_n120332# A4 a_1238_n120332# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15966 GND A4 word808 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15967 a_1370_n22636# a_1320_n66# a_1238_n22636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15968 a_710_n41096# A7 a_314_n41096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15969 a_1370_n31014# a_1320_n66# a_1238_n31014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15970 word653 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15971 GND A0 word848 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15972 GND A8 word94 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15973 word1004 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15974 GND A1 word908 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15975 word719 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15976 a_1238_n118344# A5 a_842_n118344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15977 word221 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15978 a_446_n106558# A8 a_50_n106558# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X15979 a_2162_n75460# a_2112_n66# a_2030_n75460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15980 a_1238_n109966# A5 a_974_n109966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15981 word151 a_2376_n66# a_2162_n21642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15982 a_710_n79578# A7 a_446_n79578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15983 a_1766_n61828# A3 a_1370_n61828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15984 GND A3 word1011 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15985 word1011 a_2376_n66# a_2162_n143762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15986 word817 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15987 GND A6 word23 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15988 GND A2 word155 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15989 GND A0 word746 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15990 word902 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15991 GND A8 word641 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15992 a_1370_n127006# a_1320_n66# a_1106_n127006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15993 word758 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15994 word481 a_2376_n66# a_2294_n68502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15995 GND A7 word277 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15996 GND A8 word582 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X15997 GND A1 word417 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15998 GND A8 word711 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X15999 word783 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16000 a_1766_n38966# A3 a_1370_n38966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16001 a_2294_n103576# A1 a_2030_n103576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16002 GND A2 word643 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16003 GND A1 word844 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16004 GND A3 word789 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16005 a_1238_n100878# A5 a_842_n100878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16006 word911 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16007 GND A1 word785 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16008 GND A2 word152 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16009 GND A2 word211 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16010 a_1106_n50752# a_1056_n66# a_842_n50752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16011 word789 a_2376_n66# a_2294_n112238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16012 word270 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16013 a_2030_n52598# A2 a_1766_n52598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16014 word985 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16015 a_1106_n97612# a_1056_n66# a_974_n97612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16016 word984 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16017 word428 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16018 GND A2 word482 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16019 GND A4 word972 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16020 GND A1 word353 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16021 a_2030_n99458# A2 a_1634_n99458# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16022 a_710_n123456# A7 a_314_n123456# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16023 GND A8 word38 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16024 word640 A0 a_2294_n91080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16025 GND A8 word760 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16026 GND A8 word199 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16027 GND A7 word543 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16028 a_446_n94630# A8 a_50_n94630# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16029 a_1766_n85116# A3 a_1370_n85116# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16030 GND A1 word624 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16031 word847 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16032 a_446_n33286# A8 a_182_n33286# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16033 GND A1 word192 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16034 GND A8 word687 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16035 a_446_n9004# A8 a_182_n9004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16036 word920 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16037 GND A9 word295 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16038 a_2030_n90370# A2 a_1634_n90370# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16039 GND A8 word757 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16040 a_2294_n118486# A1 a_2030_n118486# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16041 GND A5 word6 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16042 GND A7 word57 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16043 a_2162_n5028# a_2112_n66# a_2030_n5028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16044 word818 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16045 GND A3 word835 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16046 GND A2 word257 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16047 a_1370_n75318# a_1320_n66# a_1238_n75318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16048 a_710_n85400# A7 a_446_n85400# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16049 word835 a_2376_n66# a_2162_n118770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16050 a_578_n138082# a_528_n66# a_314_n138082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16051 GND A4 word747 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16052 a_1238_n342# A5 a_974_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16053 a_1370_n66940# a_1320_n66# a_1238_n66940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16054 word858 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16055 GND A5 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16056 a_974_n96902# A6 a_578_n96902# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16057 word799 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16058 word463 a_2376_n66# a_2162_n65946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16059 GND A7 word318 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16060 GND A0 word728 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16061 a_974_n7158# A6 a_710_n7158# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16062 a_50_n114936# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16063 a_50_n123314# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16064 a_1766_n53166# A3 a_1370_n53166# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16065 GND A7 word259 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16066 GND A5 word860 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16067 a_1106_n34138# a_1056_n66# a_842_n34138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16068 GND A8 word521 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16069 a_1106_n25760# a_1056_n66# a_974_n25760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16070 GND A6 word158 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16071 word952 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16072 a_182_n47912# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16073 GND A5 word916 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16074 GND A2 word523 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16075 GND A6 word646 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16076 a_1502_n141064# A4 a_1106_n141064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16077 GND A5 word857 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16078 GND A0 word160 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16079 GND A2 word722 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16080 a_1502_n132686# A4 a_1106_n132686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16081 a_710_n120900# A7 a_314_n120900# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16082 a_1370_n43368# a_1320_n66# a_1106_n43368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16083 GND A0 word994 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16084 word53 a_2376_n66# a_2294_n7726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16085 a_842_n35416# a_792_n66# a_578_n35416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16086 a_1370_n34990# a_1320_n66# a_1106_n34990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16087 GND A8 word240 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16088 GND A7 word525 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16089 GND A7 word584 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16090 a_1238_n139076# A5 a_842_n139076# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16091 word297 a_2376_n66# a_2294_n42374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16092 a_1766_n82560# A3 a_1502_n82560# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16093 GND A1 word665 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16094 word148 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16095 word946 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16096 a_314_n45924# a_264_n66# a_182_n45924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16097 a_314_n54302# a_264_n66# a_182_n54302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16098 word89 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16099 GND A0 word216 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16100 GND A1 word233 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16101 word697 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16102 GND A6 word424 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16103 word627 a_2376_n66# a_2162_n89234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16104 a_1370_n139360# a_1320_n66# a_1238_n139360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16105 a_50_n138224# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16106 word986 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16107 word927 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16108 a_446_n6448# A8 a_182_n6448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16109 a_50_n129846# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16110 GND A0 word546 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16111 word636 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16112 a_446_n77590# A8 a_50_n77590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16113 a_1766_n59698# A3 a_1502_n59698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16114 GND A5 word965 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16115 word412 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16116 a_182_n15962# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16117 word143 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16118 GND A8 word626 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16119 GND A6 word263 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16120 a_1106_n71484# a_1056_n66# a_842_n71484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16121 word800 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16122 word859 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16123 a_578_n63532# a_528_n66# a_314_n63532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16124 a_1370_n81140# a_1320_n66# a_1106_n81140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16125 word766 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16126 a_50_n85826# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16127 a_50_n94204# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16128 word57 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16129 a_842_n64810# a_792_n66# a_578_n64810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16130 word633 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16131 GND A0 word324 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16132 GND A7 word359 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16133 word563 a_2376_n66# a_2162_n80146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16134 GND A2 word827 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16135 a_50_n120758# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16136 GND A7 word300 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16137 word536 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16138 GND A1 word440 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16139 GND A4 word258 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16140 a_1370_n49900# a_1320_n66# a_1238_n49900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16141 a_1370_n58278# a_1320_n66# a_1238_n58278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16142 word61 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16143 GND A7 word630 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16144 word829 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16145 a_578_n23630# a_528_n66# a_446_n23630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16146 a_578_n32008# a_528_n66# a_446_n32008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16147 a_842_n72762# a_792_n66# a_578_n72762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16148 a_974_n79862# A6 a_710_n79862# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16149 a_842_n103718# a_792_n66# a_578_n103718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16150 a_50_n106274# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16151 word253 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16152 a_182_n53734# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16153 a_182_n62112# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16154 a_314_n69212# a_264_n66# a_182_n69212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16155 word706 A0 a_2162_n100452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16156 a_314_n115504# a_264_n66# a_50_n115504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16157 GND A6 word529 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16158 a_1106_n17098# a_1056_n66# a_842_n17098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16159 GND A4 word995 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16160 a_578_n92926# a_528_n66# a_446_n92926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16161 a_578_n31582# a_528_n66# a_446_n31582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16162 a_842_n32860# a_792_n66# a_578_n32860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16163 a_974_n39960# A6 a_710_n39960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16164 word964 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16165 word962 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16166 a_182_n4034# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16167 a_182_n22210# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16168 GND A4 word524 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16169 GND A6 word526 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16170 a_314_n51746# a_264_n66# a_182_n51746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16171 a_314_n60124# a_264_n66# a_182_n60124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16172 word928 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16173 word945 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16174 GND A3 word66 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16175 word810 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16176 a_50_n144046# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16177 word609 a_2376_n66# a_2294_n86678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16178 a_50_n135668# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16179 GND A1 word545 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16180 a_1502_n73614# A4 a_1238_n73614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16181 a_182_n30162# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16182 a_314_n37262# a_264_n66# a_182_n37262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16183 word453 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16184 word826 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16185 a_182_n21784# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16186 a_842_n87672# a_792_n66# a_710_n87672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16187 a_842_n127006# a_792_n66# a_710_n127006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16188 GND A6 word304 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16189 word866 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16190 a_842_n118628# a_792_n66# a_710_n118628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16191 a_578_n60976# a_528_n66# a_314_n60976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16192 GND A3 word262 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16193 word807 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16194 a_710_n2188# A7 a_446_n2188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16195 a_182_n68644# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16196 a_50_n91648# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16197 word455 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16198 word752 A0 a_2294_n106984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16199 a_1634_n4460# a_1584_n66# a_1370_n4460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16200 a_2294_n5880# A1 a_2030_n5880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16201 word796 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16202 word577 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16203 word737 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16204 GND A4 word358 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16205 word518 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16206 a_50_n77164# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16207 GND A4 word299 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16208 a_842_n47770# a_792_n66# a_710_n47770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16209 a_974_n94062# A6 a_578_n94062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16210 word870 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16211 GND A0 word204 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16212 word511 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16213 a_182_n37120# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16214 a_50_n112096# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16215 a_1502_n19228# A4 a_1238_n19228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16216 a_314_n66656# a_264_n66# a_182_n66656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16217 GND A4 word197 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16218 a_1106_n133112# a_1056_n66# a_974_n133112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16219 a_1106_n124734# a_1056_n66# a_842_n124734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16220 GND A4 word138 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16221 a_1502_n41664# A4 a_1106_n41664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16222 a_314_n112948# a_264_n66# a_50_n112948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16223 a_314_n121326# a_264_n66# a_50_n121326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16224 GND A6 word570 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16225 GND A0 word692 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16226 a_1502_n1336# A4 a_1238_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16227 word186 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16228 a_1502_n88524# A4 a_1106_n88524# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16229 a_2030_n8578# A2 a_1634_n8578# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16230 word1018 A0 a_2162_n144756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16231 word926 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16232 a_182_n45072# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16233 a_182_n36694# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16234 word230 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16235 GND A6 word409 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16236 a_2030_n104712# A2 a_1766_n104712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16237 word411 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16238 word1003 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16239 GND A0 word140 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16240 word971 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16241 a_182_n1478# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16242 a_1502_n10140# A4 a_1238_n10140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16243 a_1898_n57994# a_1848_n66# a_1766_n57994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16244 a_1238_n65804# A5 a_842_n65804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16245 word251 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16246 word901 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16247 a_50_n141490# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16248 word391 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16249 word623 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16250 word842 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16251 word682 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16252 GND A2 word914 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16253 word29 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16254 a_314_n43084# a_264_n66# a_182_n43084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16255 word189 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16256 word494 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16257 word435 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16258 a_1898_n133822# a_1848_n66# a_1634_n133822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16259 word130 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16260 word975 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16261 a_842_n124450# a_792_n66# a_710_n124450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16262 word340 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16263 GND A3 word244 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16264 a_1502_n56574# A4 a_1238_n56574# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16265 a_314_n136236# a_264_n66# a_50_n136236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16266 GND A6 word675 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16267 word852 A0 a_2294_n121184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16268 a_314_n127858# a_264_n66# a_50_n127858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16269 word677 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16270 word333 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16271 GND A0 word16 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16272 GND A6 word912 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16273 word778 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16274 GND A2 word850 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16275 a_2030_n119622# A2 a_1634_n119622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16276 a_974_n128710# A6 a_578_n128710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16277 word335 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16278 a_578_n99174# a_528_n66# a_446_n99174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16279 a_1634_n81424# a_1584_n66# a_1370_n81424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16280 GND A2 word34 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16281 a_1502_n25050# A4 a_1106_n25050# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16282 word298 A0 a_2162_n42516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16283 a_1106_n108120# a_1056_n66# a_842_n108120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16284 a_314_n72478# a_264_n66# a_182_n72478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16285 a_1634_n131124# a_1584_n66# a_1370_n131124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16286 word234 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16287 a_1634_n122746# a_1584_n66# a_1370_n122746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16288 a_1898_n101872# a_1848_n66# a_1634_n101872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16289 word227 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16290 a_1634_n58562# a_1584_n66# a_1370_n58562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16291 word750 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16292 word196 A0 a_2294_n28032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16293 a_1634_n108262# a_1584_n66# a_1370_n108262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16294 a_1106_n116072# a_1056_n66# a_974_n116072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16295 a_1106_n107694# a_1056_n66# a_842_n107694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16296 word452 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16297 a_842_n139360# a_792_n66# a_578_n139360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16298 a_2030_n110534# A2 a_1634_n110534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16299 a_1370_n8578# a_1320_n66# a_1106_n8578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16300 GND A5 word448 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16301 GND A3 word566 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16302 GND A9 word441 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16303 a_1238_n10282# A5 a_842_n10282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16304 a_2294_n70632# A1 a_2030_n70632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16305 a_710_n45214# A7 a_314_n45214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16306 a_1634_n27038# a_1584_n66# a_1370_n27038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16307 word351 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16308 a_710_n36836# A7 a_314_n36836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16309 GND A5 word346 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16310 word883 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16311 word664 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16312 word748 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16313 a_1238_n57142# A5 a_974_n57142# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16314 a_2162_n103434# a_2112_n66# a_1898_n103434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16315 a_1238_n48764# A5 a_842_n48764# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16316 a_1898_n108830# a_1848_n66# a_1634_n108830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16317 word622 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16318 a_2162_n18234# a_2112_n66# a_1898_n18234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16319 word493 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16320 word434 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16321 a_1634_n87956# a_1584_n66# a_1502_n87956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16322 word271 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16323 word339 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16324 a_314_n142058# a_264_n66# a_50_n142058# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16325 GND A9 word160 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16326 a_1106_n145466# a_1056_n66# a_842_n145466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16327 a_1634_n137656# a_1584_n66# a_1502_n137656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16328 word70 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16329 a_314_n133680# a_264_n66# a_50_n133680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16330 word659 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16331 a_1238_n9288# A5 a_842_n9288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16332 a_1898_n116782# a_1848_n66# a_1766_n116782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16333 GND A5 word282 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16334 GND A3 word615 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16335 GND A6 word953 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16336 GND A5 word223 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16337 GND A3 word183 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16338 GND A7 word806 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16339 a_2030_n125444# A2 a_1766_n125444# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16340 a_2294_n16246# A1 a_2030_n16246# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16341 a_710_n74608# A7 a_446_n74608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16342 a_314_n119196# a_264_n66# a_50_n119196# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16343 GND A9 word216 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16344 word639 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16345 a_2162_n132828# a_2112_n66# a_1898_n132828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16346 a_710_n13264# A7 a_446_n13264# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16347 a_2162_n47628# a_2112_n66# a_1898_n47628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16348 a_2294_n85542# A1 a_2030_n85542# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16349 GND A8 word67 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16350 word537 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16351 word610 A0 a_2162_n86820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16352 GND A4 word550 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16353 a_1502_n91790# A4 a_1238_n91790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16354 word1011 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16355 word178 A0 a_2162_n25476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16356 word114 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16357 GND A9 word324 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16358 GND A9 word265 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16359 word107 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16360 GND A3 word390 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16361 word666 A0 a_2162_n94772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16362 a_1766_n114368# A3 a_1502_n114368# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16363 a_2294_n45640# A1 a_2030_n45640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16364 a_710_n42658# A7 a_314_n42658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16365 a_2030_n33144# A2 a_1634_n33144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16366 a_710_n51036# A7 a_314_n51036# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16367 word602 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16368 GND A5 word328 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16369 GND A5 word387 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16370 word730 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16371 a_1238_n119906# A5 a_842_n119906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16372 GND A4 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16373 a_710_n89518# A7 a_446_n89518# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16374 word604 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16375 GND A9 word321 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16376 a_2294_n53592# A1 a_2030_n53592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16377 word444 A0 a_2294_n63248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16378 word913 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16379 word972 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16380 word853 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16381 a_1766_n48906# A3 a_1370_n48906# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16382 GND A8 word722 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16383 word53 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16384 word314 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16385 word373 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16386 a_1634_n79294# a_1584_n66# a_1502_n79294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16387 GND A7 word22 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16388 GND A7 word847 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16389 GND A6 word935 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16390 GND A2 word281 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16391 GND A4 word712 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16392 a_1238_n110818# A5 a_974_n110818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16393 GND A9 word99 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16394 a_2030_n131266# A2 a_1634_n131266# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16395 a_578_n133112# a_528_n66# a_314_n133112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16396 word6 A0 a_2162_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16397 a_710_n80430# A7 a_446_n80430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16398 a_2030_n122888# A2 a_1766_n122888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16399 GND A5 word594 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16400 a_1238_n83980# A5 a_842_n83980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16401 a_1238_n92358# A5 a_974_n92358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16402 a_2162_n53450# a_2112_n66# a_1898_n53450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16403 GND A1 word753 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16404 a_1502_n136804# A4 a_1238_n136804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16405 a_2030_n48054# A2 a_1766_n48054# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16406 word519 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16407 word835 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16408 word894 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16409 word396 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16410 word747 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16411 a_2162_n115788# a_2112_n66# a_1898_n115788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16412 GND A7 word122 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16413 a_2294_n142910# A1 a_1898_n142910# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16414 a_1766_n25334# A3 a_1370_n25334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16415 a_446_n34848# A8 a_182_n34848# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16416 a_1766_n16956# A3 a_1370_n16956# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16417 GND A9 word37 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16418 a_974_n1762# A6 a_710_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16419 word490 A0 a_2162_n69780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16420 GND A9 word365 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16421 word899 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16422 a_2162_n99884# a_2112_n66# a_1898_n99884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16423 a_578_n101162# a_528_n66# a_446_n101162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16424 GND A5 word17 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16425 word419 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16426 GND A7 word68 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16427 GND A2 word386 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16428 word829 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16429 GND A9 word204 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16430 GND A1 word960 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16431 word905 a_2376_n66# a_2294_n128710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16432 a_578_n139644# a_528_n66# a_314_n139644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16433 a_2162_n21500# a_2112_n66# a_1898_n21500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16434 a_2294_n28600# A1 a_2030_n28600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16435 a_2030_n77448# A2 a_1766_n77448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16436 a_1502_n104854# A4 a_1106_n104854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16437 a_2030_n137798# A2 a_1634_n137798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16438 word52 A0 a_2294_n7584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16439 word603 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16440 word954 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16441 word1013 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16442 GND A0 word798 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16443 word171 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16444 GND A7 word329 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16445 a_974_n8720# A6 a_710_n8720# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16446 word101 a_2376_n66# a_2294_n14542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16447 a_1766_n54728# A3 a_1502_n54728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16448 a_2294_n97896# A1 a_2030_n97896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16449 GND A1 word1016 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16450 GND A3 word961 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16451 a_2162_n90796# a_2112_n66# a_1898_n90796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16452 word683 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16453 word961 a_2376_n66# a_2294_n136662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16454 a_2294_n110960# A1 a_1898_n110960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16455 a_446_n11276# A8 a_182_n11276# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16456 a_1370_n84832# a_1320_n66# a_1238_n84832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16457 a_2162_n139076# a_2112_n66# a_2030_n139076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16458 word767 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16459 GND A2 word105 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16460 a_578_n108120# a_528_n66# a_446_n108120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16461 GND A8 word591 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16462 GND A8 word532 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16463 GND A9 word140 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16464 word733 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16465 word1022 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16466 word685 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16467 a_578_n130556# a_528_n66# a_314_n130556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16468 word22 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16469 a_446_n80572# A8 a_50_n80572# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16470 GND A2 word593 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16471 GND A5 word986 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16472 GND A5 word927 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16473 a_1238_n102156# A5 a_842_n102156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16474 GND A3 word739 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16475 a_1502_n142626# A4 a_1106_n142626# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16476 a_1766_n135100# A3 a_1370_n135100# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16477 GND A2 word161 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16478 a_1106_n43652# a_1056_n66# a_974_n43652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16479 word739 a_2376_n66# a_2162_n105138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16480 a_1370_n53308# a_1320_n66# a_1106_n53308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16481 a_578_n107694# a_528_n66# a_446_n107694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16482 a_1370_n44930# a_1320_n66# a_1106_n44930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16483 word703 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16484 word367 a_2376_n66# a_2162_n52314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16485 word378 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16486 a_1370_n102440# a_1320_n66# a_1238_n102440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16487 a_710_n116356# A7 a_314_n116356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16488 a_1502_n128142# A4 a_1238_n128142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16489 a_1502_n119764# A4 a_1238_n119764# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16490 a_50_n101304# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16491 GND A7 word104 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16492 GND A0 word286 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16493 GND A1 word244 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16494 GND A5 word705 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16495 GND A9 word19 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16496 word999 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16497 a_1370_n52882# a_1320_n66# a_1106_n52882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16498 a_1766_n78016# A3 a_1502_n78016# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16499 a_446_n87530# A8 a_50_n87530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16500 a_2294_n134248# A1 a_2030_n134248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16501 word797 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16502 a_710_n484# A7 a_446_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16503 a_2294_n125870# A1 a_1898_n125870# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16504 a_182_n25902# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16505 a_446_n26186# A8 a_182_n26186# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16506 GND A1 word28 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16507 a_1370_n99742# a_1320_n66# a_1106_n99742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16508 GND A8 word696 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16509 a_1106_n81424# a_1056_n66# a_974_n81424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16510 word870 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16511 word929 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16512 a_1238_n131550# A5 a_974_n131550# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16513 GND A2 word368 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16514 a_578_n145466# a_528_n66# a_314_n145466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16515 a_710_n6306# A7 a_446_n6306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16516 a_2030_n83270# A2 a_1634_n83270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16517 a_1502_n110676# A4 a_1238_n110676# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16518 a_446_n95482# A8 a_50_n95482# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16519 a_1370_n21358# a_1320_n66# a_1238_n21358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16520 GND A2 word698 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16521 word995 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16522 a_842_n13406# a_792_n66# a_710_n13406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16523 a_1370_n12980# a_1320_n66# a_1238_n12980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16524 GND A8 word85 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16525 GND A7 word370 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16526 word768 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16527 GND A1 word840 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16528 GND A0 word780 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16529 a_974_n42942# A6 a_710_n42942# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16530 a_446_n105280# A8 a_50_n105280# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16531 word83 a_2376_n66# a_2162_n11986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16532 a_710_n78300# A7 a_446_n78300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16533 a_1370_n68218# a_1320_n66# a_1238_n68218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16534 word926 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16535 GND A6 word14 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16536 word542 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16537 a_1370_n90654# a_1320_n66# a_1106_n90654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16538 a_842_n82702# a_792_n66# a_710_n82702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16539 GND A8 word573 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16540 a_1370_n117350# a_1320_n66# a_1106_n117350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16541 a_50_n116214# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16542 word413 a_2376_n66# a_2294_n58846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16543 GND A7 word268 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16544 word1004 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16545 a_50_n107836# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16546 a_1766_n46066# A3 a_1502_n46066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16547 GND A1 word349 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16548 GND A1 word408 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16549 GND A2 word634 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16550 a_1106_n27038# a_1056_n66# a_974_n27038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16551 a_1370_n67792# a_1320_n66# a_1238_n67792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16552 a_974_n80714# A6 a_710_n80714# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16553 a_1106_n96334# a_1056_n66# a_974_n96334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16554 word975 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16555 GND A0 word110 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16556 GND A2 word473 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16557 a_1106_n87956# a_1056_n66# a_842_n87956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16558 a_2030_n98180# A2 a_1766_n98180# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16559 GND A2 word731 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16560 GND A4 word904 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16561 a_710_n122178# A7 a_314_n122178# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16562 a_710_n113800# A7 a_314_n113800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16563 word998 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16564 GND A4 word162 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16565 GND A1 word285 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16566 word1015 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16567 GND A4 word103 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16568 a_842_n28316# a_792_n66# a_578_n28316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16569 a_1370_n36268# a_1320_n66# a_1106_n36268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16570 GND A8 word190 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16571 word679 a_2376_n66# a_2162_n96618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16572 GND A7 word534 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16573 GND A0 word944 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16574 a_974_n57852# A6 a_578_n57852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16575 a_2030_n3608# A2 a_1634_n3608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16576 word247 a_2376_n66# a_2162_n35274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16577 a_842_n50752# a_792_n66# a_710_n50752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16578 a_1766_n75460# A3 a_1370_n75460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16579 a_2294_n140070# A1 a_2030_n140070# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16580 a_314_n47202# a_264_n66# a_182_n47202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16581 word1 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16582 GND A0 word166 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16583 a_182_n31724# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16584 a_314_n38824# a_264_n66# a_182_n38824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16585 a_182_n40102# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16586 a_1502_n13832# A4 a_1106_n13832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16587 GND A6 word315 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16588 GND A8 word678 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16589 a_4348_164# A5 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X16590 a_1898_n61402# a_1848_n66# a_1634_n61402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16591 a_578_n70916# a_528_n66# a_314_n70916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16592 a_710_n3750# A7 a_446_n3750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16593 word822 A0 a_2162_n116924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16594 word93 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16595 a_974_n26328# A6 a_578_n26328# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16596 a_842_n10850# a_792_n66# a_710_n10850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16597 GND A2 word680 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16598 word809 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16599 a_578_n56432# a_528_n66# a_314_n56432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16600 a_50_n87104# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16601 a_50_n78726# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16602 word790 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16603 GND A0 word274 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16604 word513 a_2376_n66# a_2294_n73046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16605 word581 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16606 a_974_n95624# A6 a_578_n95624# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16607 GND A5 word971 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16608 VDD A2 a_1848_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X16609 a_50_n122036# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16610 a_1898_n4318# a_1848_n66# a_1634_n4318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16611 word305 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16612 GND A7 word309 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16613 GND A6 word701 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16614 a_50_n113658# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16615 GND A0 word432 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16616 GND A4 word267 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16617 a_1502_n51604# A4 a_1106_n51604# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16618 word298 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16619 GND A6 word149 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16620 a_842_n65662# a_792_n66# a_578_n65662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16621 word151 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16622 word711 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16623 word996 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16624 a_182_n55012# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16625 a_182_n46634# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16626 a_1502_n28742# A4 a_1238_n28742# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16627 GND A6 word420 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16628 word481 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16629 GND A0 word210 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16630 a_1898_n67934# a_1848_n66# a_1634_n67934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16631 a_578_n94204# a_528_n66# a_446_n94204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16632 GND A2 word514 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16633 GND A2 word713 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16634 word691 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16635 word982 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16636 word632 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16637 a_578_n24482# a_528_n66# a_446_n24482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16638 a_842_n34138# a_792_n66# a_578_n34138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16639 word198 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16640 a_1766_n5028# A3 a_1502_n5028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16641 a_974_n63674# A6 a_578_n63674# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16642 a_1106_n79294# a_1056_n66# a_974_n79294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16643 word912 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16644 GND A2 word984 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16645 word774 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16646 word356 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16647 word693 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16648 GND A9 a_0_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X16649 a_182_n15110# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16650 a_314_n53024# a_264_n66# a_182_n53024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16651 word80 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16652 word937 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16653 word878 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16654 a_314_n44646# a_264_n66# a_182_n44646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16655 word686 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16656 word505 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16657 word895 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16658 GND A4 word47 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16659 a_1898_n36410# a_1848_n66# a_1634_n36410# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16660 word559 a_2376_n66# a_2162_n79578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16661 a_1370_n3608# a_1320_n66# a_1238_n3608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16662 a_50_n128568# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16663 word410 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16664 word918 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16665 a_446_n5170# A8 a_182_n5170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16666 word568 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16667 word922 A0 a_2162_n131124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16668 word403 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16669 a_182_n23062# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16670 a_182_n14684# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16671 word848 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16672 GND A2 word920 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16673 a_578_n62254# a_528_n66# a_314_n62254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16674 a_842_n142342# a_792_n66# a_578_n142342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16675 a_1898_n35984# a_1848_n66# a_1634_n35984# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16676 a_1898_n44362# a_1848_n66# a_1766_n44362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16677 word466 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16678 a_974_n79010# A6 a_710_n79010# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16679 a_50_n84548# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16680 word405 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16681 word407 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16682 a_2294_n7158# A1 a_2030_n7158# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16683 GND A2 word619 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16684 word96 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16685 word495 a_2376_n66# a_2162_n70490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16686 word746 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16687 GND A2 word818 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16688 word527 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16689 a_5140_164# A8 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X16690 a_842_n49048# a_792_n66# a_710_n49048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16691 word879 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16692 a_1238_n4318# A5 a_974_n4318# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16693 a_842_n71484# a_792_n66# a_578_n71484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16694 word461 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16695 a_974_n78584# A6 a_710_n78584# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16696 word820 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16697 a_842_n102440# a_792_n66# a_578_n102440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16698 a_1502_n95908# A4 a_1106_n95908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16699 GND A3 word148 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16700 word185 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16701 a_1106_n126012# a_1056_n66# a_842_n126012# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16702 a_182_n52456# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16703 a_314_n59556# a_264_n66# a_182_n59556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16704 a_314_n114226# a_264_n66# a_50_n114226# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16705 GND A6 word520 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16706 a_1634_n118202# a_1584_n66# a_1370_n118202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16707 a_1106_n117634# a_1056_n66# a_974_n117634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16708 word463 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16709 a_1898_n73756# a_1848_n66# a_1766_n73756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16710 a_578_n91648# a_528_n66# a_446_n91648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16711 word1023 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16712 GND A5 word86 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16713 word968 A0 a_2294_n137656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16714 word876 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16715 a_1238_n3892# A5 a_974_n3892# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16716 a_1238_n20222# A5 a_974_n20222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16717 a_182_n29594# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16718 a_1238_n11844# A5 a_842_n11844# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16719 word239 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16720 word362 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16721 word631 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16722 word180 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16723 word953 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16724 GND A4 word515 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16725 a_50_n99458# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16726 a_578_n68786# a_528_n66# a_314_n68786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16727 a_1238_n58704# A5 a_974_n58704# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16728 a_314_n50468# a_264_n66# a_182_n50468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16729 word79 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16730 a_842_n17098# a_792_n66# a_710_n17098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16731 a_50_n134390# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16732 word201 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16733 GND A0 word578 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16734 a_974_n114652# A6 a_710_n114652# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16735 word341 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16736 GND A3 word355 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16737 a_1502_n63958# A4 a_1238_n63958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16738 a_314_n143620# a_264_n66# a_50_n143620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16739 word444 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16740 word47 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16741 word567 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16742 word385 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16743 GND A6 word295 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16744 a_842_n86394# a_792_n66# a_710_n86394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16745 a_1898_n19370# a_1848_n66# a_1766_n19370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16746 word238 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16747 GND A3 word194 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16748 word507 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16749 word802 A0 a_2162_n114084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16750 a_182_n58988# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16751 a_182_n67366# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16752 a_50_n90370# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16753 a_314_n129136# a_264_n66# a_50_n129136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16754 GND A9 word286 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16755 a_2162_n10708# a_2112_n66# a_2030_n10708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16756 a_2294_n17808# A1 a_1898_n17808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16757 a_710_n14826# A7 a_446_n14826# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16758 word406 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16759 a_1898_n88666# a_1848_n66# a_1634_n88666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16760 GND A2 word859 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16761 GND A2 word800 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16762 GND A5 word132 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16763 word728 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16764 GND A4 word290 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16765 word467 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16766 word502 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16767 a_1634_n74324# a_1584_n66# a_1502_n74324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16768 a_1634_n65946# a_1584_n66# a_1502_n65946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16769 GND A4 word620 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16770 a_2162_n119906# a_2112_n66# a_2030_n119906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16771 a_182_n9288# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16772 word248 A0 a_2294_n35416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16773 a_314_n57000# a_264_n66# a_182_n57000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16774 a_314_n65378# a_264_n66# a_182_n65378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16775 a_314_n120048# a_264_n66# a_50_n120048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16776 a_1634_n124024# a_1584_n66# a_1502_n124024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16777 a_1106_n123456# a_1056_n66# a_842_n123456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16778 a_1634_n115646# a_1584_n66# a_1502_n115646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16779 a_314_n111670# a_264_n66# a_50_n111670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16780 word504 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16781 a_974_n129562# A6 a_578_n129562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16782 a_2030_n7300# A2 a_1766_n7300# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16783 word118 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16784 word177 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16785 a_1502_n87246# A4 a_1106_n87246# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16786 GND A6 word798 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16787 a_1502_n78868# A4 a_1106_n78868# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16788 GND A4 word676 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16789 word490 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16790 a_2030_n34706# A2 a_1766_n34706# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16791 word402 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16792 word935 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16793 word994 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16794 GND A5 word398 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16795 a_2162_n110818# a_2112_n66# a_2030_n110818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16796 a_1238_n64526# A5 a_842_n64526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16797 word712 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16798 a_2162_n25618# a_2112_n66# a_2030_n25618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16799 GND A3 word516 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16800 GND A9 word391 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16801 word119 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16802 a_710_n38114# A7 a_314_n38114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16803 word242 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16804 word833 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16805 a_1766_n123882# A3 a_1502_n123882# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16806 a_1634_n33996# a_1584_n66# a_1502_n33996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16807 a_1634_n42374# a_1584_n66# a_1502_n42374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16808 word614 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16809 word20 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16810 GND A4 word395 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16811 word856 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16812 a_2162_n94914# a_2112_n66# a_2030_n94914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16813 a_1898_n132544# a_1848_n66# a_1766_n132544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16814 word443 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16815 word607 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16816 GND A9 word110 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16817 a_2030_n141206# A2 a_1766_n141206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16818 a_2294_n23630# A1 a_1898_n23630# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16819 a_2294_n32008# A1 a_2030_n32008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16820 a_1502_n55296# A4 a_1238_n55296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16821 a_314_n126580# a_264_n66# a_50_n126580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16822 word668 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16823 word447 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16824 word506 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16825 a_1502_n6590# A4 a_1106_n6590# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16826 a_1238_n93920# A5 a_974_n93920# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16827 GND A6 word903 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16828 a_1766_n139218# A3 a_1370_n139218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16829 GND A3 word133 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16830 a_1898_n101020# a_1848_n66# a_1766_n101020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16831 a_1106_n5312# a_1056_n66# a_974_n5312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16832 GND A2 word131 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16833 word508 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16834 a_2294_n92926# A1 a_1898_n92926# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16835 a_2030_n118344# A2 a_1766_n118344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16836 word589 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16837 word449 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16838 GND A9 word166 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16839 a_2162_n134106# a_2112_n66# a_1898_n134106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16840 a_2294_n31582# A1 a_1898_n31582# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16841 a_1634_n71768# a_1584_n66# a_1370_n71768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16842 word157 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16843 word230 A0 a_2162_n32860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16844 word758 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16845 a_314_n71200# a_264_n66# a_182_n71200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16846 word347 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16847 a_1766_n138792# A3 a_1370_n138792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16848 a_974_n135384# A6 a_578_n135384# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16849 a_2162_n62964# a_2112_n66# a_2030_n62964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16850 word487 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16851 word560 A0 a_2294_n79720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16852 word555 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16853 a_1502_n93068# A4 a_1238_n93068# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16854 GND A6 word780 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16855 word128 A0 a_2294_n18376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16856 word961 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16857 a_1766_n130130# A3 a_1370_n130130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16858 a_578_n102724# a_528_n66# a_446_n102724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16859 word489 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16860 word548 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16861 a_1370_n7300# a_1320_n66# a_1106_n7300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16862 GND A9 word274 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16863 GND A3 word340 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16864 word616 A0 a_2294_n87672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16865 a_1766_n107268# A3 a_1370_n107268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16866 GND A9 word432 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16867 a_2030_n17666# A2 a_1634_n17666# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16868 GND A5 word337 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16869 word423 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16870 a_2294_n60976# A1 a_1898_n60976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16871 GND A5 word278 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16872 a_2162_n102156# a_2112_n66# a_1898_n102156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16873 word739 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16874 a_1238_n47486# A5 a_842_n47486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16875 word613 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16876 GND A9 word271 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16877 a_446_n21216# A8 a_182_n21216# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16878 GND A6 word43 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16879 a_1634_n95056# a_1584_n66# a_1370_n95056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16880 a_446_n12838# A8 a_182_n12838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16881 word394 A0 a_2162_n56148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16882 word425 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16883 a_2030_n86962# A2 a_1766_n86962# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16884 GND A9 word210 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16885 word803 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16886 word330 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16887 GND A8 word731 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16888 a_1370_n143904# a_1320_n66# a_1106_n143904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16889 a_1106_n144188# a_1056_n66# a_842_n144188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16890 a_1634_n136378# a_1584_n66# a_1370_n136378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16891 a_446_n90512# A8 a_50_n90512# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16892 GND A8 word111 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16893 a_2162_n77874# a_2112_n66# a_2030_n77874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16894 a_2162_n86252# a_2112_n66# a_1898_n86252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16895 a_2294_n106416# A1 a_1898_n106416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16896 word650 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16897 a_446_n108972# A8 a_50_n108972# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16898 GND A5 word214 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16899 GND A6 word944 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16900 GND A1 word805 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16901 a_446_n100310# A8 a_50_n100310# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16902 a_1238_n103718# A5 a_842_n103718# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16903 GND A7 word797 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16904 a_710_n73330# A7 a_446_n73330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16905 a_2030_n124166# A2 a_1634_n124166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16906 a_1238_n85258# A5 a_842_n85258# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16907 a_1238_n76880# A5 a_974_n76880# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16908 GND A5 word836 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16909 a_710_n117918# A7 a_314_n117918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16910 a_1766_n32718# A3 a_1502_n32718# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16911 GND A8 word58 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16912 a_2294_n75886# A1 a_1898_n75886# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16913 a_2294_n84264# A1 a_2030_n84264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16914 GND A1 word861 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16915 GND A3 word806 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16916 word346 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16917 a_710_n81282# A7 a_446_n81282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16918 a_1370_n62822# a_1320_n66# a_1106_n62822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16919 word469 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16920 a_2162_n117066# a_2112_n66# a_1898_n117066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16921 word1002 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16922 word808 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16923 a_1370_n111954# a_1320_n66# a_1238_n111954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16924 a_446_n27748# A8 a_182_n27748# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16925 a_446_n36126# A8 a_182_n36126# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16926 a_710_n41380# A7 a_314_n41380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16927 word282 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16928 GND A8 word155 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16929 word223 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16930 a_1106_n68502# a_1056_n66# a_842_n68502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16931 a_2030_n139076# A2 a_1766_n139076# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16932 a_1238_n118628# A5 a_842_n118628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16933 word153 a_2376_n66# a_2294_n21926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16934 a_710_n88240# A7 a_446_n88240# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16935 a_1502_n106132# A4 a_1106_n106132# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16936 word595 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16937 word996 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16938 GND A1 word148 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16939 a_1634_n92500# a_1584_n66# a_1502_n92500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16940 GND A1 word89 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16941 GND A6 word25 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16942 word553 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16943 GND A0 word748 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16944 GND A8 word643 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16945 word904 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16946 word121 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16947 a_1370_n30872# a_1320_n66# a_1238_n30872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16948 GND A8 word211 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16949 GND A7 word279 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16950 a_2294_n99174# A1 a_2030_n99174# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16951 GND A8 word713 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16952 a_1634_n142200# a_1584_n66# a_1502_n142200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16953 word785 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16954 a_2162_n7442# a_2112_n66# a_2030_n7442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16955 GND A8 word152 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16956 GND A1 word636 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16957 a_2162_n92074# a_2112_n66# a_1898_n92074# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16958 a_2294_n112238# A1 a_1898_n112238# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16959 word911 a_2376_n66# a_2162_n129562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16960 GND A7 word13 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16961 GND A8 word541 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16962 word774 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16963 word972 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16964 a_1370_n135242# a_1320_n66# a_1106_n135242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16965 a_1370_n126864# a_1320_n66# a_1106_n126864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16966 GND A5 word585 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16967 a_446_n73472# A8 a_50_n73472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16968 a_1238_n91080# A5 a_974_n91080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16969 GND A4 word974 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16970 a_710_n123740# A7 a_314_n123740# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16971 a_974_n20932# A6 a_578_n20932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16972 a_2294_n90086# A1 a_2030_n90086# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16973 GND A8 word40 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16974 word847 a_2376_n66# a_2162_n120474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16975 word317 a_2376_n66# a_2294_n45214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16976 word328 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16977 GND A7 word113 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16978 a_710_n109256# A7 a_314_n109256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16979 a_446_n33570# A8 a_182_n33570# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16980 GND A0 word236 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16981 GND A1 word253 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16982 GND A9 word28 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16983 GND A7 word601 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16984 GND A8 word759 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16985 a_1766_n93352# A3 a_1370_n93352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16986 a_1370_n103292# a_1320_n66# a_1238_n103292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16987 word747 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16988 a_446_n19086# A8 a_182_n19086# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16989 a_1766_n84974# A3 a_1370_n84974# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X16990 a_182_n18802# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16991 GND A5 word8 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16992 GND A7 word59 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16993 word879 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16994 word820 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16995 GND A5 word711 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16996 GND A2 word259 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16997 GND A6 word441 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X16998 a_578_n138366# a_528_n66# a_314_n138366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X16999 a_578_n129988# a_528_n66# a_314_n129988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17000 GND A4 word749 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17001 a_1238_n626# A5 a_974_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17002 word860 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17003 a_446_n8862# A8 a_182_n8862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17004 GND A5 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17005 a_446_n88382# A8 a_50_n88382# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17006 GND A5 word982 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17007 GND A4 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17008 GND A7 word379 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17009 GND A0 word730 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17010 word945 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17011 GND A1 word460 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17012 GND A7 word320 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17013 a_1766_n53450# A3 a_1370_n53450# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17014 word876 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17015 word741 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17016 GND A6 word160 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17017 GND A8 word523 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17018 word916 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17019 word857 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17020 a_50_n109114# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17021 word722 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17022 word954 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17023 GND A7 word376 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17024 word64 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17025 GND A1 word516 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17026 GND A2 word584 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17027 a_1502_n141348# A4 a_1106_n141348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17028 GND A5 word918 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17029 a_1502_n132970# A4 a_1106_n132970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17030 a_578_n34422# a_528_n66# a_446_n34422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17031 a_1106_n33996# a_1056_n66# a_842_n33996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17032 a_1106_n42374# a_1056_n66# a_974_n42374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17033 a_1238_n139360# A5 a_842_n139360# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17034 a_974_n73614# A6 a_710_n73614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17035 a_1106_n89234# a_1056_n66# a_842_n89234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17036 GND A6 word546 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17037 a_50_n100026# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17038 GND A7 word95 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17039 word299 a_2376_n66# a_2162_n42658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17040 a_710_n115078# A7 a_314_n115078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17041 a_1502_n118486# A4 a_1238_n118486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17042 a_1766_n21500# A3 a_1370_n21500# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17043 word948 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17044 word699 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17045 GND A0 word894 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17046 word629 a_2376_n66# a_2294_n89518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17047 a_50_n138508# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17048 word197 a_2376_n66# a_2294_n28174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17049 a_1766_n68360# A3 a_1502_n68360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17050 GND A7 word583 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17051 a_182_n33002# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17052 GND A0 word116 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17053 GND A1 word133 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17054 a_1370_n98464# a_1320_n66# a_1106_n98464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17055 a_182_n24624# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17056 word1021 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17057 GND A8 word628 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17058 GND A6 word265 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17059 a_1106_n71768# a_1056_n66# a_842_n71768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17060 a_1106_n80146# a_1056_n66# a_974_n80146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17061 word886 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17062 a_578_n63816# a_528_n66# a_314_n63816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17063 a_1898_n54302# a_1848_n66# a_1634_n54302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17064 word536 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17065 a_842_n143904# a_792_n66# a_578_n143904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17066 word827 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17067 a_578_n144188# a_528_n66# a_314_n144188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17068 a_710_n5028# A7 a_446_n5028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17069 word32 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17070 word477 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17071 GND A1 word621 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17072 word772 A0 a_2294_n109824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17073 GND A3 word22 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17074 word59 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17075 word635 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17076 GND A2 word689 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17077 a_842_n12128# a_792_n66# a_710_n12128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17078 a_2294_n8720# A1 a_1898_n8720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17079 a_974_n19228# A6 a_578_n19228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17080 word565 a_2376_n66# a_2294_n80430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17081 a_974_n41664# A6 a_710_n41664# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17082 a_1370_n80998# a_1320_n66# a_1106_n80998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17083 GND A8 word564 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17084 a_50_n106558# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17085 word255 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17086 GND A0 word382 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17087 a_1634_n6874# a_1584_n66# a_1502_n6874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17088 GND A1 word340 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17089 word708 A0 a_2294_n100736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17090 a_1898_n22352# a_1848_n66# a_1634_n22352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17091 a_842_n120332# a_792_n66# a_710_n120332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17092 a_578_n31866# a_528_n66# a_446_n31866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17093 a_182_n39534# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17094 word311 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17095 word252 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17096 GND A2 word464 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17097 a_1898_n69212# a_1848_n66# a_1766_n69212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17098 a_1106_n86678# a_1056_n66# a_842_n86678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17099 a_182_n4318# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17100 a_314_n60408# a_264_n66# a_182_n60408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17101 word81 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17102 GND A3 word68 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17103 GND A0 word648 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17104 word724 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17105 a_50_n144330# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17106 a_974_n56574# A6 a_578_n56574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17107 word887 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17108 GND A4 word582 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17109 GND A4 word641 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17110 word455 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17111 word828 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17112 a_182_n3892# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17113 a_182_n30446# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17114 a_314_n37546# a_264_n66# a_182_n37546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17115 GND A8 word669 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17116 a_1898_n29310# a_1848_n66# a_1634_n29310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17117 a_842_n87956# a_792_n66# a_710_n87956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17118 word146 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17119 a_1898_n60124# a_1848_n66# a_1766_n60124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17120 word872 A0 a_2294_n124024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17121 a_182_n68928# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17122 a_1502_n59414# A4 a_1106_n59414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17123 GND A0 word36 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17124 word46 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17125 word84 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17126 a_974_n25050# A6 a_578_n25050# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17127 GND A4 word421 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17128 a_1898_n98606# a_1848_n66# a_1766_n98606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17129 word511 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17130 GND A2 word929 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17131 word206 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17132 word579 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17133 word798 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17134 a_1898_n37262# a_1848_n66# a_1766_n37262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17135 a_578_n55154# a_528_n66# a_314_n55154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17136 GND A4 word360 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17137 a_842_n126864# a_792_n66# a_710_n126864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17138 a_50_n77448# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17139 a_974_n94346# A6 a_578_n94346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17140 word572 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17141 word445 a_2376_n66# a_2294_n63390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17142 GND A2 word768 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17143 GND A6 word692 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17144 a_50_n112380# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17145 a_1898_n3040# a_1848_n66# a_1766_n3040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17146 a_314_n66940# a_264_n66# a_182_n66940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17147 a_1502_n50326# A4 a_1106_n50326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17148 GND A0 word364 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17149 GND A4 word199 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17150 a_1502_n41948# A4 a_1106_n41948# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17151 a_314_n121610# a_264_n66# a_50_n121610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17152 word576 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17153 word289 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17154 GND A4 word357 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17155 a_1502_n1620# A4 a_1238_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17156 GND A6 word140 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17157 a_842_n64384# a_792_n66# a_578_n64384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17158 word142 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17159 GND A0 word694 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17160 a_182_n45356# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17161 GND A3 word98 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17162 GND A4 word687 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17163 a_182_n36978# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17164 GND A2 word51 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17165 a_1502_n27464# A4 a_1238_n27464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17166 word472 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17167 word251 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17168 a_1898_n75034# a_1848_n66# a_1634_n75034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17169 word413 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17170 word1005 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17171 a_1898_n66656# a_1848_n66# a_1766_n66656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17172 GND A6 word569 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17173 GND A2 word704 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17174 word914 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17175 a_842_n103292# a_792_n66# a_578_n103292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17176 a_1238_n13122# A5 a_842_n13122# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17177 word35 a_2376_n66# a_2162_n5170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17178 word189 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17179 word903 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17180 a_974_n130414# A6 a_578_n130414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17181 a_1634_n52314# a_1584_n66# a_1502_n52314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17182 a_974_n62396# A6 a_578_n62396# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17183 word684 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17184 word625 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17185 a_314_n43368# a_264_n66# a_182_n43368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17186 a_1634_n102014# a_1584_n66# a_1502_n102014# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17187 word869 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17188 word677 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17189 GND A4 word38 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17190 a_50_n127290# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17191 a_1634_n29452# a_1584_n66# a_1502_n29452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17192 GND A0 word528 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17193 word850 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17194 GND A3 word305 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17195 a_1502_n56858# A4 a_1238_n56858# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17196 a_1502_n65236# A4 a_1238_n65236# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17197 a_314_n136520# a_264_n66# a_50_n136520# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17198 word854 A0 a_2162_n121468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17199 GND A4 word521 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17200 word679 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17201 word394 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17202 word335 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17203 GND A0 word18 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17204 word247 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17205 word780 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17206 a_1898_n43084# a_1848_n66# a_1634_n43084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17207 word188 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17208 a_842_n141064# a_792_n66# a_578_n141064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17209 a_50_n83270# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17210 GND A9 word236 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17211 a_2030_n119906# A2 a_1634_n119906# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17212 a_710_n16104# A7 a_446_n16104# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17213 a_578_n99458# a_528_n66# a_446_n99458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17214 a_314_n144472# a_264_n66# a_50_n144472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17215 a_1634_n81708# a_1584_n66# a_1370_n81708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17216 a_974_n91790# A6 a_578_n91790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17217 GND A2 word809 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17218 word227 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17219 word87 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17220 a_1634_n20364# a_1584_n66# a_1502_n20364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17221 a_1238_n28032# A5 a_842_n28032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17222 GND A3 word691 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17223 a_1634_n131408# a_1584_n66# a_1370_n131408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17224 a_1238_n19654# A5 a_974_n19654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17225 a_1238_n3040# A5 a_974_n3040# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17226 word229 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17227 a_1634_n58846# a_1584_n66# a_1370_n58846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17228 word452 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17229 a_1634_n67224# a_1584_n66# a_1370_n67224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17230 word198 A0 a_2162_n28316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17231 a_182_n51178# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17232 a_314_n58278# a_264_n66# a_182_n58278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17233 GND A3 word80 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17234 a_1106_n116356# a_1056_n66# a_974_n116356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17235 a_3556_164# A2 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X17236 a_182_n42800# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17237 a_314_n49900# a_264_n66# a_182_n49900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17238 GND A2 word33 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17239 word134 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17240 a_1502_n33286# A4 a_1106_n33286# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17241 word356 A0 a_2294_n50752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17242 a_1106_n107978# a_1056_n66# a_842_n107978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17243 a_1634_n108546# a_1584_n66# a_1370_n108546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17244 a_2030_n110818# A2 a_1634_n110818# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17245 word351 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17246 word454 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17247 word1014 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17248 a_1634_n130982# a_1584_n66# a_1370_n130982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17249 GND A5 word77 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17250 word127 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17251 a_1898_n72478# a_1848_n66# a_1634_n72478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17252 word686 A0 a_2162_n97612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17253 word664 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17254 word900 A0 a_2294_n128000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17255 a_1238_n10566# A5 a_842_n10566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17256 word622 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17257 a_2030_n27606# A2 a_1766_n27606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17258 word353 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17259 word944 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17260 GND A5 word348 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17261 word493 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17262 word885 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17263 a_1238_n57426# A5 a_974_n57426# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17264 a_50_n98180# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17265 word624 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17266 GND A9 word341 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17267 word70 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17268 GND A3 word407 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17269 GND A3 word466 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17270 a_2162_n40954# a_2112_n66# a_1898_n40954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17271 word192 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17272 a_2294_n56432# A1 a_1898_n56432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17273 a_2030_n96902# A2 a_1634_n96902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17274 a_974_n113374# A6 a_710_n113374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17275 a_1766_n116782# A3 a_1370_n116782# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17276 a_1634_n26896# a_1584_n66# a_1370_n26896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17277 word273 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17278 word38 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17279 GND A8 word181 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17280 a_1634_n137940# a_1584_n66# a_1502_n137940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17281 word557 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17282 GND A5 word284 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17283 GND A6 word955 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17284 GND A7 word867 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17285 a_182_n66088# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17286 GND A7 word808 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17287 a_314_n119480# a_264_n66# a_50_n119480# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17288 a_710_n13548# A7 a_446_n13548# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17289 a_1898_n87388# a_1848_n66# a_1766_n87388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17290 word719 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17291 GND A3 word673 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17292 word458 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17293 GND A9 word116 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17294 a_2030_n64952# A2 a_1634_n64952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17295 a_710_n82844# A7 a_446_n82844# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17296 word539 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17297 word767 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17298 a_2162_n118628# a_2112_n66# a_2030_n118628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17299 a_314_n64100# a_264_n66# a_182_n64100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17300 word107 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17301 word180 A0 a_2294_n25760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17302 a_1238_n94772# A5 a_974_n94772# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17303 word175 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17304 a_2162_n64242# a_2112_n66# a_2030_n64242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17305 a_1634_n105990# a_1584_n66# a_1502_n105990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17306 a_1106_n113800# a_1056_n66# a_974_n113800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17307 word495 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17308 a_974_n128284# A6 a_578_n128284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17309 a_974_n4602# A6 a_710_n4602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17310 word168 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17311 GND A6 word789 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17312 word109 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17313 a_1502_n77590# A4 a_1106_n77590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17314 word1000 A0 a_2294_n142200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17315 a_1766_n123030# A3 a_1502_n123030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17316 a_578_n104002# a_528_n66# a_446_n104002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17317 word663 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17318 a_2030_n33428# A2 a_1634_n33428# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17319 a_710_n51320# A7 a_314_n51320# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17320 word985 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17321 GND A5 word389 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17322 word703 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17323 a_1238_n54870# A5 a_974_n54870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17324 GND A9 word382 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17325 a_2162_n24340# a_2112_n66# a_2030_n24340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17326 word233 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17327 a_2294_n62254# A1 a_1898_n62254# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17328 word373 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17329 word974 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17330 a_4348_164# A5 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X17331 word191 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17332 a_1370_n40812# a_1320_n66# a_1238_n40812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17333 a_710_n50894# A7 a_314_n50894# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17334 word855 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17335 GND A8 word222 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17336 a_2162_n93636# a_2112_n66# a_2030_n93636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17337 word712 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17338 word847 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17339 GND A3 word981 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17340 GND A1 word977 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17341 word981 a_2376_n66# a_2294_n139502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17342 a_446_n14116# A8 a_182_n14116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17343 a_2162_n32292# a_2112_n66# a_2030_n32292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17344 a_2294_n39392# A1 a_1898_n39392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17345 word375 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17346 a_1634_n79578# a_1584_n66# a_1502_n79578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17347 a_2030_n79862# A2 a_1766_n79862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17348 GND A7 word24 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17349 word344 A0 a_2294_n49048# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17350 word502 A0 a_2162_n71484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17351 word753 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17352 GND A7 word849 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17353 a_1634_n129278# a_1584_n66# a_1502_n129278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17354 GND A5 word655 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17355 word8 A0 a_2294_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17356 a_446_n83412# A8 a_50_n83412# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17357 word438 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17358 a_2294_n121752# A1 a_2030_n121752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17359 GND A2 word122 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17360 a_1238_n31298# A5 a_842_n31298# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17361 word499 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17362 a_2294_n91648# A1 a_1898_n91648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17363 GND A3 word917 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17364 a_2030_n48338# A2 a_1766_n48338# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17365 GND A9 word157 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17366 word917 a_2376_n66# a_2294_n130414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17367 a_2030_n39960# A2 a_1634_n39960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17368 a_1634_n70490# a_1584_n66# a_1502_n70490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17369 a_2030_n70774# A2 a_1766_n70774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17370 word398 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17371 GND A5 word652 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17372 a_2162_n124450# a_2112_n66# a_2030_n124450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17373 word702 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17374 word749 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17375 GND A9 word487 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17376 GND A7 word124 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17377 a_2162_n39250# a_2112_n66# a_2030_n39250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17378 a_1634_n120190# a_1584_n66# a_1502_n120190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17379 a_1766_n25618# A3 a_1370_n25618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17380 word338 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17381 a_446_n101162# A8 a_50_n101162# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17382 GND A1 word752 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17383 GND A3 word756 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17384 a_710_n74182# A7 a_446_n74182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17385 word419 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17386 GND A9 word39 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17387 a_2294_n128710# A1 a_2030_n128710# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17388 a_1370_n113232# a_1320_n66# a_1238_n113232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17389 a_446_n29026# A8 a_182_n29026# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17390 a_578_n101446# a_528_n66# a_446_n101446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17391 GND A1 word48 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17392 word480 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17393 word638 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17394 GND A5 word781 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17395 GND A2 word329 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17396 GND A9 word423 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17397 GND A5 word722 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17398 VDD A9 a_0_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X17399 a_710_n110108# A7 a_314_n110108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17400 GND A9 word364 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17401 a_578_n139928# a_528_n66# a_314_n139928# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17402 word54 A0 a_2162_n7868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17403 a_1106_n14542# a_1056_n66# a_842_n14542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17404 a_446_n89944# A8 a_50_n89944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17405 a_446_n98322# A8 a_50_n98322# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17406 a_2030_n16388# A2 a_1766_n16388# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17407 GND A5 word269 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17408 word1015 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17409 a_2294_n136662# A1 a_2030_n136662# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17410 word232 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17411 GND A8 word105 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17412 a_446_n108120# A8 a_50_n108120# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17413 word173 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17414 word946 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17415 GND A3 word963 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17416 word103 a_2376_n66# a_2162_n14826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17417 a_446_n11560# A8 a_182_n11560# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17418 GND A6 word34 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17419 a_1634_n85400# a_1584_n66# a_1370_n85400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17420 a_2030_n85684# A2 a_1634_n85684# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17421 word685 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17422 word963 a_2376_n66# a_2162_n136946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17423 word986 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17424 GND A8 word593 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17425 word927 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17426 GND A0 word856 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17427 GND A8 word102 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17428 GND A8 word161 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17429 word735 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17430 a_578_n130840# a_528_n66# a_314_n130840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17431 a_1766_n71342# A3 a_1370_n71342# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17432 a_446_n107694# A8 a_50_n107694# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17433 a_2162_n76596# a_2112_n66# a_2030_n76596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17434 word24 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17435 a_446_n80856# A8 a_50_n80856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17436 a_710_n89092# A7 a_446_n89092# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17437 a_1502_n142910# A4 a_1106_n142910# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17438 GND A2 word163 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17439 a_1106_n43936# a_1056_n66# a_974_n43936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17440 a_1106_n52314# a_1056_n66# a_842_n52314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17441 a_1238_n102440# A5 a_842_n102440# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17442 GND A7 word788 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17443 word766 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17444 GND A2 word104 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17445 GND A6 word286 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17446 a_578_n107978# a_528_n66# a_446_n107978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17447 GND A5 word535 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17448 a_1502_n128426# A4 a_1238_n128426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17449 a_710_n125018# A7 a_314_n125018# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17450 a_1634_n1904# a_1584_n66# a_1502_n1904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17451 GND A1 word305 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17452 a_710_n116640# A7 a_314_n116640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17453 GND A2 word651 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17454 GND A9 word469 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17455 GND A1 word852 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17456 a_1370_n39108# a_1320_n66# a_1238_n39108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17457 a_710_n49190# A7 a_314_n49190# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17458 GND A8 word49 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17459 a_1238_n110392# A5 a_974_n110392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17460 GND A3 word738 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17461 word797 a_2376_n66# a_2294_n113374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17462 a_1370_n61544# a_1320_n66# a_1106_n61544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17463 word267 a_2376_n66# a_2162_n38114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17464 word858 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17465 a_710_n768# A7 a_446_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17466 GND A0 word186 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17467 word799 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17468 a_446_n26470# A8 a_182_n26470# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17469 a_710_n124592# A7 a_314_n124592# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17470 GND A1 word361 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17471 GND A8 word698 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17472 GND A2 word370 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17473 a_1106_n81708# a_1056_n66# a_974_n81708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17474 GND A8 word207 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17475 GND A7 word551 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17476 a_1502_n110960# A4 a_1238_n110960# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17477 a_446_n95766# A8 a_50_n95766# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17478 a_1766_n77874# A3 a_1502_n77874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17479 GND A1 word632 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17480 a_1370_n30020# a_1320_n66# a_1238_n30020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17481 word770 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17482 GND A6 word391 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17483 word987 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17484 GND A2 word209 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17485 word928 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17486 GND A1 word80 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17487 GND A2 word426 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17488 a_1370_n90938# a_1320_n66# a_1106_n90938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17489 GND A8 word634 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17490 GND A7 word270 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17491 GND A8 word575 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17492 a_1766_n46350# A3 a_1502_n46350# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17493 GND A8 word704 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17494 GND A1 word957 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17495 GND A3 word902 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17496 word35 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17497 a_2162_n6164# a_2112_n66# a_2030_n6164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17498 GND A1 word568 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17499 word826 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17500 a_1370_n76454# a_1320_n66# a_1238_n76454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17501 a_842_n68502# a_792_n66# a_578_n68502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17502 word731 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17503 word904 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17504 GND A2 word145 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17505 a_1898_n23914# a_1848_n66# a_1766_n23914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17506 word381 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17507 GND A7 word326 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17508 a_1370_n125586# a_1320_n66# a_1106_n125586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17509 a_446_n1052# A8 a_182_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17510 a_1898_n6732# a_1848_n66# a_1634_n6732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17511 a_974_n8294# A6 a_710_n8294# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17512 a_1106_n96618# a_1056_n66# a_974_n96618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17513 GND A2 word475 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17514 GND A4 word965 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17515 a_1106_n35274# a_1056_n66# a_842_n35274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17516 a_578_n18944# a_528_n66# a_446_n18944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17517 a_578_n27322# a_528_n66# a_446_n27322# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17518 a_1106_n26896# a_1056_n66# a_974_n26896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17519 GND A6 word166 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17520 word319 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17521 word249 a_2376_n66# a_2294_n35558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17522 word3 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17523 a_1766_n14400# A3 a_1502_n14400# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17524 GND A1 word185 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17525 GND A4 word67 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17526 GND A8 word680 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17527 a_446_n8010# A8 a_182_n8010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17528 GND A0 word1002 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17529 word61 a_2376_n66# a_2294_n8862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17530 GND A7 word533 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17531 GND A7 word592 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17532 GND A8 word750 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17533 word791 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17534 a_1766_n7442# A3 a_1370_n7442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17535 a_1766_n92074# A3 a_1502_n92074# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17536 GND A1 word673 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17537 a_182_n17524# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17538 word156 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17539 GND A4 word491 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17540 GND A7 word50 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17541 GND A6 word274 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17542 GND A6 word432 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17543 a_842_n136804# a_792_n66# a_578_n136804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17544 a_578_n137088# a_528_n66# a_314_n137088# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17545 GND A4 word740 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17546 word41 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17547 GND A2 word250 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17548 a_578_n56716# a_528_n66# a_314_n56716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17549 a_1502_n102298# A4 a_1238_n102298# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17550 a_446_n7584# A8 a_182_n7584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17551 word585 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17552 word515 a_2376_n66# a_2162_n73330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17553 a_974_n95908# A6 a_578_n95908# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17554 GND A5 word973 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17555 a_50_n122320# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17556 GND A5 word914 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17557 word151 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17558 GND A0 word434 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17559 GND A6 word271 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17560 word646 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17561 GND A4 word427 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17562 a_50_n86962# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17563 word212 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17564 GND A8 word514 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17565 a_842_n65946# a_792_n66# a_578_n65946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17566 word153 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17567 word998 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17568 a_1634_n8152# a_1584_n66# a_1370_n8152# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17569 GND A0 word332 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17570 word571 a_2376_n66# a_2162_n81282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17571 a_182_n46918# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17572 a_50_n121894# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17573 a_50_n130272# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17574 a_1502_n37404# A4 a_1238_n37404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17575 GND A4 word266 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17576 GND A2 word715 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17577 word356 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17578 GND A5 word850 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17579 a_1106_n41096# a_1056_n66# a_974_n41096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17580 word693 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17581 a_578_n24766# a_528_n66# a_446_n24766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17582 a_578_n33144# a_528_n66# a_446_n33144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17583 a_842_n104854# a_792_n66# a_578_n104854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17584 word8 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17585 a_1106_n79578# a_1056_n66# a_974_n79578# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17586 GND A6 word537 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17587 word939 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17588 a_314_n44930# a_264_n66# a_182_n44930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17589 a_314_n53308# a_264_n66# a_182_n53308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17590 a_50_n137230# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17591 GND A0 word598 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17592 a_842_n33996# a_792_n66# a_578_n33996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17593 GND A7 word633 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17594 word924 A0 a_2294_n131408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17595 a_1766_n4886# A3 a_1502_n4886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17596 word67 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17597 GND A4 word591 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17598 a_182_n23346# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17599 word405 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17600 a_182_n14968# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17601 a_842_n89234# a_792_n66# a_710_n89234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17602 GND A8 word619 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17603 a_314_n52882# a_264_n66# a_182_n52882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17604 a_1898_n53024# a_1848_n66# a_1766_n53024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17605 a_1106_n70490# a_1056_n66# a_842_n70490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17606 a_842_n142626# a_792_n66# a_578_n142626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17607 word818 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17608 a_50_n93210# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17609 a_50_n145182# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17610 a_578_n62538# a_528_n66# a_314_n62538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17611 word759 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17612 word468 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17613 word50 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17614 word748 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17615 word461 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17616 a_1766_n111812# A3 a_1370_n111812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17617 a_974_n40386# A6 a_710_n40386# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17618 word529 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17619 a_1634_n21926# a_1584_n66# a_1370_n21926# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17620 a_842_n119764# a_792_n66# a_710_n119764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17621 a_50_n92784# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17622 word463 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17623 a_974_n78868# A6 a_710_n78868# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17624 a_842_n71768# a_792_n66# a_578_n71768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17625 word395 a_2376_n66# a_2162_n56290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17626 a_314_n68218# a_264_n66# a_182_n68218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17627 a_50_n105280# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17628 GND A0 word314 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17629 a_182_n52740# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17630 a_314_n59840# a_264_n66# a_182_n59840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17631 a_182_n61118# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17632 a_1502_n43226# A4 a_1106_n43226# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17633 a_314_n114510# a_264_n66# a_50_n114510# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17634 a_1106_n117918# a_1056_n66# a_974_n117918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17635 GND A4 word366 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17636 word526 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17637 a_1634_n140922# a_1584_n66# a_1370_n140922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17638 word362 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17639 word970 A0 a_2162_n137940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17640 word878 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17641 a_578_n30588# a_528_n66# a_446_n30588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17642 a_1238_n20506# A5 a_974_n20506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17643 a_182_n38256# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17644 a_182_n29878# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17645 a_182_n60692# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17646 a_314_n67792# a_264_n66# a_182_n67792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17647 word955 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17648 GND A9 word81 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17649 a_314_n122462# a_264_n66# a_50_n122462# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17650 a_182_n3040# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17651 GND A6 word519 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17652 a_974_n55296# A6 a_578_n55296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17653 a_974_n114936# A6 a_710_n114936# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17654 word238 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17655 a_1634_n45214# a_1584_n66# a_1370_n45214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17656 word343 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17657 GND A0 word580 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17658 word1011 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17659 word819 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17660 a_1502_n11276# A4 a_1238_n11276# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17661 a_182_n20790# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17662 a_842_n86678# a_792_n66# a_710_n86678# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17663 GND A0 word478 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17664 word859 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17665 word509 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17666 a_182_n67650# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17667 a_314_n129420# a_264_n66# a_50_n129420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17668 word344 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17669 word804 A0 a_2294_n114368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17670 word37 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17671 word467 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17672 a_1502_n9430# A4 a_1238_n9430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17673 word197 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17674 a_1898_n97328# a_1848_n66# a_1634_n97328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17675 word789 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17676 word502 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17677 GND A5 word193 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17678 word138 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17679 word570 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17680 word730 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17681 word983 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17682 a_1370_n3182# a_1320_n66# a_1238_n3182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17683 a_842_n125586# a_792_n66# a_710_n125586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17684 a_50_n76170# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17685 GND A3 word311 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17686 GND A9 word186 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17687 a_2294_n34422# A1 a_2030_n34422# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17688 a_1634_n74608# a_1584_n66# a_1502_n74608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17689 a_314_n137372# a_264_n66# a_50_n137372# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17690 a_974_n93068# A6 a_578_n93068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17691 a_314_n128994# a_264_n66# a_50_n128994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17692 GND A6 word683 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17693 a_1634_n13264# a_1584_n66# a_1370_n13264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17694 word177 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17695 a_1106_n132118# a_1056_n66# a_974_n132118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17696 a_1634_n124308# a_1584_n66# a_1502_n124308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17697 a_1106_n123740# a_1056_n66# a_842_n123740# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17698 a_2162_n65804# a_2112_n66# a_1898_n65804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17699 a_1898_n103434# a_1848_n66# a_1766_n103434# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17700 a_1634_n115930# a_1584_n66# a_1502_n115930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17701 a_974_n129846# A6 a_578_n129846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17702 word179 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17703 a_1502_n87530# A4 a_1106_n87530# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17704 word919 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17705 word981 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17706 a_182_n44078# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17707 GND A2 word42 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17708 word306 A0 a_2162_n43652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17709 word674 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17710 GND A4 word678 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17711 a_2030_n103718# A2 a_1634_n103718# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17712 a_182_n35700# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17713 word404 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17714 word242 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17715 a_1238_n64810# A5 a_842_n64810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17716 GND A3 word518 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17717 GND A3 word577 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17718 a_2294_n63816# A1 a_2030_n63816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17719 a_1766_n132544# A3 a_1502_n132544# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17720 word244 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17721 word443 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17722 word894 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17723 word835 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17724 a_1634_n42658# a_1584_n66# a_1502_n42658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17725 word675 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17726 word84 A0 a_2294_n12128# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17727 GND A5 word456 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17728 a_314_n42090# a_264_n66# a_182_n42090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17729 GND A3 word416 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17730 word668 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17731 a_1898_n132828# a_1848_n66# a_1766_n132828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17732 a_974_n99600# A6 a_578_n99600# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17733 a_1766_n109682# A3 a_1502_n109682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17734 a_1634_n19796# a_1584_n66# a_1502_n19796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17735 a_710_n37972# A7 a_314_n37972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17736 a_1502_n55580# A4 a_1238_n55580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17737 word572 A0 a_2294_n81424# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17738 a_1766_n101020# A3 a_1502_n101020# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17739 word756 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17740 GND A8 word131 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17741 word670 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17742 a_1898_n109966# a_1848_n66# a_1766_n109966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17743 word501 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17744 GND A6 word905 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17745 word442 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17746 GND A7 word817 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17747 GND A3 word135 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17748 GND A3 word352 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17749 word510 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17750 GND A9 word227 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17751 a_2030_n118628# A2 a_1766_n118628# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17752 a_314_n143194# a_264_n66# a_50_n143194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17753 word78 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17754 word347 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17755 a_578_n98180# a_528_n66# a_446_n98180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17756 a_1766_n100594# A3 a_1502_n100594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17757 a_1238_n18376# A5 a_974_n18376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17758 word159 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17759 a_2294_n87104# A1 a_1898_n87104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17760 GND A1 word881 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17761 a_2162_n71626# a_2112_n66# a_1898_n71626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17762 a_2294_n78726# A1 a_2030_n78726# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17763 a_2162_n80004# a_2112_n66# a_2030_n80004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17764 word489 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17765 word349 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17766 a_710_n84122# A7 a_446_n84122# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17767 a_446_n102724# A8 a_50_n102724# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17768 a_1898_n100878# a_1848_n66# a_1766_n100878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17769 a_974_n135668# A6 a_578_n135668# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17770 a_2162_n10282# a_2112_n66# a_1898_n10282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17771 a_2294_n17382# A1 a_2030_n17382# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17772 a_710_n75744# A7 a_446_n75744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17773 word963 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17774 word1022 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17775 word130 A0 a_2162_n18660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17776 a_2162_n133964# a_2112_n66# a_1898_n133964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17777 a_1106_n115078# a_1056_n66# a_974_n115078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17778 a_1106_n106700# a_1056_n66# a_842_n106700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17779 word445 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17780 word283 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17781 a_2162_n48764# a_2112_n66# a_1898_n48764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17782 a_1898_n71200# a_1848_n66# a_1766_n71200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17783 GND A9 word493 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17784 word950 A0 a_2162_n135100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17785 word618 A0 a_2162_n87956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17786 GND A9 word434 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17787 word554 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17788 a_710_n44220# A7 a_314_n44220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17789 a_2030_n26328# A2 a_1634_n26328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17790 GND A5 word280 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17791 GND A5 word339 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17792 word425 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17793 a_1238_n47770# A5 a_842_n47770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17794 a_1238_n56148# A5 a_974_n56148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17795 word547 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17796 word615 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17797 GND A9 word332 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17798 a_1634_n95340# a_1584_n66# a_1370_n95340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17799 a_2030_n95624# A2 a_1766_n95624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17800 GND A9 word273 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17801 a_2294_n46776# A1 a_2030_n46776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17802 a_974_n112096# A6 a_710_n112096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17803 a_710_n52172# A7 a_314_n52172# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17804 word323 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17805 GND A8 word11 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17806 a_710_n43794# A7 a_314_n43794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17807 GND A8 word231 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17808 a_1634_n145040# a_1584_n66# a_1370_n145040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17809 word805 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17810 GND A8 word172 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17811 word738 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17812 a_1766_n72904# A3 a_1502_n72904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17813 a_1898_n115788# a_1848_n66# a_1634_n115788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17814 GND A7 word799 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17815 GND A7 word858 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17816 word452 A0 a_2294_n64384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17817 a_1370_n129704# a_1320_n66# a_1238_n129704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17818 a_2030_n124450# A2 a_1634_n124450# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17819 GND A5 word605 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17820 word861 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17821 a_710_n12270# A7 a_446_n12270# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17822 a_446_n76312# A8 a_50_n76312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17823 word61 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17824 word77 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17825 GND A8 word60 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17826 word791 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17827 GND A3 word867 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17828 a_1238_n120332# A5 a_842_n120332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17829 a_2030_n72052# A2 a_1634_n72052# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17830 GND A9 word107 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17831 word867 a_2376_n66# a_2162_n123314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17832 a_1238_n111954# A5 a_974_n111954# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17833 word348 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17834 a_710_n81566# A7 a_446_n81566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17835 a_1634_n63390# a_1584_n66# a_1370_n63390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17836 GND A5 word661 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17837 GND A5 word602 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17838 word1004 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17839 a_1238_n93494# A5 a_974_n93494# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17840 word916 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17841 a_1370_n120616# a_1320_n66# a_1238_n120616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17842 a_1634_n113090# a_1584_n66# a_1370_n113090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17843 a_446_n36410# A8 a_182_n36410# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17844 a_1766_n18518# A3 a_1502_n18518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17845 GND A7 word291 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17846 GND A1 word761 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17847 a_974_n3324# A6 a_710_n3324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17848 a_2162_n54586# a_2112_n66# a_1898_n54586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17849 GND A9 word48 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17850 word100 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17851 a_1370_n48622# a_1320_n66# a_1238_n48622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17852 word595 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17853 word654 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17854 word767 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17855 a_2030_n32150# A2 a_1766_n32150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17856 a_446_n35984# A8 a_182_n35984# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17857 word284 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17858 GND A5 word731 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17859 a_2030_n79010# A2 a_1634_n79010# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17860 a_1502_n106416# A4 a_1106_n106416# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17861 word998 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17862 GND A9 word373 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17863 GND A9 word314 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17864 GND A2 word496 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17865 word907 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17866 a_2294_n52598# A1 a_2030_n52598# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17867 word965 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17868 word123 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17869 GND A8 word715 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17870 GND A8 word213 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17871 a_2162_n83980# a_2112_n66# a_1898_n83980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17872 word703 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17873 word896 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17874 GND A1 word968 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17875 GND A3 word913 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17876 word913 a_2376_n66# a_2294_n129846# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17877 GND A7 word15 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17878 a_2030_n78584# A2 a_1634_n78584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17879 GND A8 word543 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17880 word974 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17881 a_1370_n16672# a_1320_n66# a_1106_n16672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17882 GND A4 word705 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17883 word1021 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17884 a_1370_n135526# a_1320_n66# a_1106_n135526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17885 GND A0 word806 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17886 a_578_n132118# a_528_n66# a_314_n132118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17887 GND A1 word536 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17888 a_446_n2614# A8 a_182_n2614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17889 a_446_n73756# A8 a_50_n73756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17890 a_446_n82134# A8 a_50_n82134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17891 a_1766_n64242# A3 a_1502_n64242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17892 GND A1 word477 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17893 a_1106_n45214# a_1056_n66# a_974_n45214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17894 GND A2 word113 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17895 GND A3 word849 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17896 a_2030_n47060# A2 a_1634_n47060# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17897 word849 a_2376_n66# a_2294_n120758# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17898 a_578_n131692# a_528_n66# a_314_n131692# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17899 word740 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17900 GND A9 word478 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17901 GND A7 word115 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17902 GND A2 word601 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17903 a_710_n109540# A7 a_314_n109540# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17904 GND A9 word419 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17905 a_1238_n103292# A5 a_842_n103292# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17906 word747 a_2376_n66# a_2162_n106274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17907 GND A9 word30 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17908 a_1370_n54444# a_1320_n66# a_1106_n54444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17909 GND A7 word603 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17910 a_2162_n98890# a_2112_n66# a_1898_n98890# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17911 a_1370_n103576# a_1320_n66# a_1238_n103576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17912 word749 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17913 a_446_n19370# A8 a_182_n19370# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17914 GND A0 word136 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17915 a_578_n100168# a_528_n66# a_446_n100168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17916 a_1766_n93636# A3 a_1370_n93636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17917 GND A5 word10 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17918 a_1766_n32292# A3 a_1502_n32292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17919 a_710_n117492# A7 a_314_n117492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17920 GND A1 word252 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17921 GND A2 word379 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17922 word982 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17923 GND A5 word713 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17924 GND A2 word320 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17925 GND A4 word810 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17926 a_578_n138650# a_528_n66# a_314_n138650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17927 a_1238_n910# A5 a_974_n910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17928 a_446_n97044# A8 a_50_n97044# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17929 word1007 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17930 a_446_n88666# A8 a_50_n88666# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17931 word655 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17932 a_2294_n135384# A1 a_2030_n135384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17933 GND A5 word5 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17934 GND A5 word984 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17935 a_974_n44504# A6 a_710_n44504# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17936 GND A3 word1013 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17937 word878 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17938 word937 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17939 GND A1 word1009 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17940 GND A0 word72 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17941 GND A2 word376 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17942 word1013 a_2376_n66# a_2294_n144046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17943 GND A4 word866 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17944 GND A4 word807 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17945 word743 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17946 a_710_n7442# A7 a_446_n7442# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17947 a_50_n96902# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17948 GND A8 word584 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17949 word760 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17950 word652 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17951 GND A8 word525 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17952 word918 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17953 a_1370_n22494# a_1320_n66# a_1238_n22494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17954 word641 a_2376_n66# a_2294_n91222# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17955 a_842_n14542# a_792_n66# a_710_n14542# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17956 a_50_n131834# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17957 a_50_n140212# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17958 a_1766_n39250# A3 a_1370_n39250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17959 GND A7 word378 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17960 GND A1 word577 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17961 a_1766_n61686# A3 a_1370_n61686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17962 GND A5 word920 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17963 a_1106_n51036# a_1056_n66# a_842_n51036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17964 word816 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17965 word757 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17966 GND A2 word154 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17967 a_1106_n42658# a_1056_n66# a_974_n42658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17968 a_578_n34706# a_528_n66# a_446_n34706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17969 a_1898_n16814# a_1848_n66# a_1766_n16814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17970 word272 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17971 word421 a_2376_n66# a_2294_n59982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17972 GND A7 word276 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17973 a_578_n106700# a_528_n66# a_446_n106700# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17974 a_50_n108972# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17975 GND A1 word416 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17976 word430 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17977 a_1106_n89518# a_1056_n66# a_842_n89518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17978 a_50_n100310# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17979 GND A2 word642 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17980 a_1502_n118770# A4 a_1238_n118770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17981 a_2030_n342# A2 a_1766_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17982 GND A3 word788 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17983 a_3556_164# A2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X17984 a_842_n52314# a_792_n66# a_710_n52314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17985 word269 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17986 a_974_n59414# A6 a_578_n59414# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X17987 word199 a_2376_n66# a_2162_n28458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17988 word983 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17989 GND A4 word971 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17990 GND A0 word118 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17991 word357 a_2376_n66# a_2294_n50894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17992 a_182_n6732# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17993 a_182_n24908# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17994 GND A1 word352 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17995 a_1370_n98748# a_1320_n66# a_1106_n98748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X17996 GND A8 word689 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17997 a_314_n62822# a_264_n66# a_182_n62822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17998 a_1106_n80430# a_1056_n66# a_974_n80430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X17999 word1023 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18000 GND A8 word630 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18001 GND A4 word111 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18002 a_842_n29452# a_792_n66# a_578_n29452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18003 word687 a_2376_n66# a_2162_n97754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18004 GND A7 word542 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18005 GND A0 word952 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18006 word741 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18007 a_2030_n4744# A2 a_1766_n4744# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18008 a_446_n94488# A8 a_50_n94488# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18009 GND A2 word200 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18010 a_974_n41948# A6 a_710_n41948# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18011 word919 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18012 GND A3 word995 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18013 word995 a_2376_n66# a_2162_n141490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18014 a_710_n4886# A7 a_446_n4886# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18015 word465 a_2376_n66# a_2294_n66230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18016 a_50_n115220# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18017 a_842_n11986# a_792_n66# a_710_n11986# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18018 word101 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18019 GND A0 word384 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18020 GND A2 word688 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18021 GND A2 word946 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18022 word596 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18023 a_1370_n66798# a_1320_n66# a_1238_n66798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18024 a_1370_n75176# a_1320_n66# a_1238_n75176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18025 a_50_n79862# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18026 a_842_n67224# a_792_n66# a_578_n67224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18027 word162 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18028 word521 a_2376_n66# a_2294_n74182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18029 word948 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18030 word895 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18031 a_842_n120616# a_792_n66# a_710_n120616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18032 a_50_n123172# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18033 a_1898_n5454# a_1848_n66# a_1766_n5454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18034 a_1898_n22636# a_1848_n66# a_1634_n22636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18035 word313 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18036 word372 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18037 a_182_n39818# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18038 a_50_n114794# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18039 GND A1 word457 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18040 a_182_n70632# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18041 a_314_n132402# a_264_n66# a_50_n132402# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18042 GND A6 word648 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18043 GND A5 word859 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18044 word306 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18045 a_578_n26044# a_528_n66# a_446_n26044# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18046 a_1898_n91932# a_1848_n66# a_1766_n91932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18047 a_842_n106132# a_792_n66# a_578_n106132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18048 GND A6 word157 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18049 word55 a_2376_n66# a_2162_n8010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18050 word308 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18051 a_974_n56858# A6 a_578_n56858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18052 word367 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18053 a_314_n46208# a_264_n66# a_182_n46208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18054 GND A0 word218 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18055 GND A4 word643 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18056 GND A2 word721 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18057 word889 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18058 a_182_n30730# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18059 a_314_n37830# a_264_n66# a_182_n37830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18060 a_842_n35274# a_792_n66# a_578_n35274# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18061 word206 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18062 GND A0 word548 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18063 word870 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18064 word874 A0 a_2162_n124308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18065 word782 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18066 GND A4 word482 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18067 GND A1 word664 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18068 word701 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18069 a_182_n16246# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18070 word88 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18071 word147 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18072 a_314_n45782# a_264_n66# a_182_n45782# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18073 a_1106_n63390# a_1056_n66# a_974_n63390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18074 word208 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18075 a_1898_n37546# a_1848_n66# a_1766_n37546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18076 a_578_n55438# a_528_n66# a_314_n55438# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18077 GND A6 word423 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18078 a_50_n86110# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18079 a_50_n138082# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18080 word926 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18081 GND A3 word322 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18082 GND A5 word964 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18083 a_314_n138934# a_264_n66# a_50_n138934# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18084 a_974_n94630# A6 a_578_n94630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18085 word574 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18086 a_1766_n104712# A3 a_1502_n104712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18087 word411 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18088 GND A6 word694 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18089 word142 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18090 GND A2 word987 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18091 GND A2 word770 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18092 GND A4 word260 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18093 word856 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18094 GND A2 word928 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18095 word63 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18096 a_1502_n50610# A4 a_1106_n50610# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18097 word637 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18098 a_50_n94062# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18099 a_50_n85684# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18100 word345 a_2376_n66# a_2294_n49190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18101 a_842_n64668# a_792_n66# a_578_n64668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18102 word413 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18103 a_2294_n8294# A1 a_2030_n8294# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18104 word144 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18105 word989 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18106 a_182_n54018# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18107 GND A0 word264 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18108 GND A2 word826 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18109 a_182_n45640# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18110 a_1502_n27748# A4 a_1238_n27748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18111 word474 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18112 GND A4 word257 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18113 a_578_n93210# a_528_n66# a_446_n93210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18114 word975 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18115 a_1106_n141632# a_1056_n66# a_842_n141632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18116 a_1634_n133822# a_1584_n66# a_1502_n133822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18117 a_1898_n66940# a_1848_n66# a_1766_n66940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18118 word887 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18119 word625 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18120 word828 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18121 a_578_n23488# a_528_n66# a_446_n23488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18122 a_1238_n13406# A5 a_842_n13406# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18123 a_842_n103576# a_792_n66# a_578_n103576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18124 a_182_n53592# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18125 GND A3 word97 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18126 a_974_n62680# A6 a_578_n62680# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18127 a_1106_n78300# a_1056_n66# a_974_n78300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18128 a_314_n115362# a_264_n66# a_50_n115362# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18129 GND A6 word528 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18130 word905 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18131 a_314_n52030# a_264_n66# a_182_n52030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18132 GND A3 word486 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18133 a_578_n92784# a_528_n66# a_446_n92784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18134 a_1238_n82702# A5 a_842_n82702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18135 word930 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18136 a_1898_n74892# a_1848_n66# a_1634_n74892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18137 word679 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18138 word976 A0 a_2294_n138792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18139 GND A4 word40 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18140 a_974_n116214# A6 a_710_n116214# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18141 word247 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18142 a_1634_n38114# a_1584_n66# a_1502_n38114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18143 GND A0 word530 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18144 word188 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18145 a_710_n47912# A7 a_314_n47912# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18146 a_1502_n65520# A4 a_1238_n65520# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18147 word961 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18148 word58 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18149 GND A4 word523 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18150 a_182_n13690# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18151 a_182_n22068# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18152 word249 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18153 word87 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18154 a_578_n61260# a_528_n66# a_314_n61260# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18155 a_1634_n101872# a_1584_n66# a_1502_n101872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18156 word750 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18157 a_842_n141348# a_792_n66# a_578_n141348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18158 a_1898_n34990# a_1848_n66# a_1766_n34990# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18159 word754 A0 a_2162_n107268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18160 GND A3 word422 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18161 word400 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18162 a_1502_n73472# A4 a_1238_n73472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18163 a_2294_n41806# A1 a_1898_n41806# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18164 a_314_n144756# a_264_n66# a_50_n144756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18165 word452 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18166 word89 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18167 word520 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18168 word739 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18169 a_2030_n20932# A2 a_1766_n20932# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18170 word229 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18171 GND A3 word693 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18172 a_842_n118486# a_792_n66# a_710_n118486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18173 a_1238_n19938# A5 a_974_n19938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18174 a_1238_n28316# A5 a_842_n28316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18175 word45 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18176 GND A3 word261 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18177 GND A9 word136 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18178 a_842_n70490# a_792_n66# a_578_n70490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18179 word454 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18180 a_1634_n67508# a_1584_n66# a_1370_n67508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18181 a_974_n77590# A6 a_710_n77590# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18182 word636 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18183 a_2162_n11844# a_2112_n66# a_2030_n11844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18184 word127 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18185 a_2294_n18944# A1 a_1898_n18944# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18186 a_710_n15962# A7 a_446_n15962# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18187 a_1106_n125018# a_1056_n66# a_842_n125018# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18188 a_1634_n117208# a_1584_n66# a_1370_n117208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18189 a_1502_n33570# A4 a_1106_n33570# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18190 a_1634_n108830# a_1584_n66# a_1370_n108830# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18191 a_1106_n116640# a_1056_n66# a_974_n116640# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18192 word294 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18193 word1020 A0 a_2294_n145040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18194 a_1238_n2898# A5 a_974_n2898# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18195 GND A5 word79 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18196 word869 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18197 a_182_n28600# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18198 a_1238_n10850# A5 a_842_n10850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18199 a_1502_n19086# A4 a_1238_n19086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18200 word256 A0 a_2294_n36552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18201 word355 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18202 GND A9 word72 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18203 a_314_n121184# a_264_n66# a_50_n121184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18204 a_1106_n124592# a_1056_n66# a_842_n124592# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18205 word617 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18206 a_1898_n49900# a_1848_n66# a_1634_n49900# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18207 a_1238_n57710# A5 a_974_n57710# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18208 a_1502_n1194# A4 a_1238_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18209 GND A3 word50 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18210 GND A3 word468 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18211 a_1502_n88382# A4 a_1106_n88382# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18212 GND A9 word343 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18213 GND A6 word806 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18214 GND A5 word76 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18215 word253 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18216 a_974_n113658# A6 a_710_n113658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18217 a_1766_n125444# A3 a_1370_n125444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18218 word194 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18219 word393 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18220 a_1634_n35558# a_1584_n66# a_1370_n35558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18221 a_2030_n35842# A2 a_1634_n35842# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18222 a_710_n53734# A7 a_314_n53734# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18223 word867 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18224 word1002 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18225 GND A5 word406 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18226 a_1898_n134106# a_1848_n66# a_1634_n134106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18227 a_2162_n120332# a_2112_n66# a_1898_n120332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18228 a_2162_n111954# a_2112_n66# a_2030_n111954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18229 a_1238_n65662# A5 a_842_n65662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18230 a_1898_n125728# a_1848_n66# a_1766_n125728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18231 a_2162_n26754# a_2112_n66# a_2030_n26754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18232 a_2162_n35132# a_2112_n66# a_1898_n35132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18233 a_842_n85400# a_792_n66# a_710_n85400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18234 word559 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18235 word522 A0 a_2162_n74324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18236 word500 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18237 word931 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18238 word28 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18239 word399 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18240 word458 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18241 word460 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18242 GND A9 word177 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18243 GND A9 word118 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18244 a_2030_n142342# A2 a_1634_n142342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18245 a_2294_n33144# A1 a_2030_n33144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18246 word495 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18247 a_314_n136094# a_264_n66# a_50_n136094# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18248 word676 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18249 a_2294_n24766# A1 a_1898_n24766# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18250 word109 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18251 word986 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18252 a_1370_n11702# a_1320_n66# a_1238_n11702# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18253 GND A6 word911 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18254 word927 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18255 a_446_n104002# A8 a_50_n104002# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18256 a_1898_n102156# a_1848_n66# a_1634_n102156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18257 a_974_n128568# A6 a_578_n128568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18258 GND A1 word772 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18259 a_710_n77022# A7 a_446_n77022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18260 word170 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18261 a_1634_n81282# a_1584_n66# a_1370_n81282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18262 word597 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18263 word972 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18264 a_2162_n135242# a_2112_n66# a_1898_n135242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18265 a_2030_n102440# A2 a_1766_n102440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18266 word766 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18267 word238 A0 a_2162_n33996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18268 word395 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18269 word705 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18270 GND A9 word443 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18271 word226 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18272 GND A9 word384 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18273 word977 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18274 GND A0 word64 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18275 a_710_n37120# A7 a_314_n37120# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18276 word235 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18277 GND A1 word708 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18278 a_2294_n139502# A1 a_1898_n139502# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18279 a_1766_n122888# A3 a_1502_n122888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18280 word375 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18281 a_2030_n110392# A2 a_1634_n110392# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18282 a_1238_n49048# A5 a_842_n49048# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18283 word556 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18284 word849 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18285 a_1238_n136804# A5 a_842_n136804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18286 a_1898_n131550# a_1848_n66# a_1634_n131550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18287 a_2294_n48054# A1 a_2030_n48054# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18288 a_1634_n88240# a_1584_n66# a_1502_n88240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18289 a_710_n112522# A7 a_314_n112522# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18290 GND A4 word836 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18291 a_710_n45072# A7 a_314_n45072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18292 a_710_n36694# A7 a_314_n36694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18293 a_1370_n26612# a_1320_n66# a_1106_n26612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18294 word681 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18295 word755 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18296 word504 A0 a_2294_n71768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18297 GND A8 word122 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18298 a_2162_n79436# a_2112_n66# a_1898_n79436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18299 a_2162_n103292# a_2112_n66# a_1898_n103292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18300 word747 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18301 word10 A0 a_2162_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18302 word499 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18303 a_1898_n108688# a_1848_n66# a_1634_n108688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18304 a_1898_n117066# a_1848_n66# a_1766_n117066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18305 a_2162_n18092# a_2112_n66# a_1898_n18092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18306 word621 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18307 a_2294_n130414# A1 a_1898_n130414# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18308 a_446_n22352# A8 a_182_n22352# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18309 GND A6 word51 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18310 word492 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18311 a_446_n13974# A8 a_182_n13974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18312 word433 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18313 word402 A0 a_2162_n57284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18314 GND A9 word218 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18315 GND A9 word159 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18316 a_2030_n117350# A2 a_1634_n117350# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18317 word811 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18318 word338 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18319 a_578_n141632# a_528_n66# a_314_n141632# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18320 a_2294_n107552# A1 a_1898_n107552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18321 GND A3 word614 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18322 GND A9 word489 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18323 a_2294_n77448# A1 a_2030_n77448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18324 GND A6 word952 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18325 GND A1 word872 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18326 GND A3 word817 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18327 a_2162_n61970# a_2112_n66# a_2030_n61970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18328 a_2162_n70348# a_2112_n66# a_1898_n70348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18329 word340 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18330 a_446_n101446# A8 a_50_n101446# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18331 a_974_n134390# A6 a_578_n134390# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18332 word817 a_2376_n66# a_2294_n116214# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18333 GND A1 word813 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18334 a_1238_n113232# A5 a_974_n113232# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18335 GND A3 word758 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18336 a_1634_n56290# a_1584_n66# a_1502_n56290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18337 a_710_n74466# A7 a_446_n74466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18338 word1013 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18339 word456 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18340 a_1238_n86394# A5 a_842_n86394# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18341 word722 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18342 a_578_n101730# a_528_n66# a_446_n101730# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18343 a_1370_n113516# a_1320_n66# a_1238_n113516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18344 a_446_n29310# A8 a_182_n29310# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18345 GND A1 word381 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18346 GND A8 word66 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18347 word668 A0 a_2294_n95056# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18348 a_1106_n23204# a_1056_n66# a_974_n23204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18349 GND A9 word425 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18350 a_1106_n14826# a_1056_n66# a_842_n14826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18351 a_446_n98606# A8 a_50_n98606# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18352 GND A5 word330 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18353 a_446_n28884# A8 a_182_n28884# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18354 word234 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18355 GND A9 word323 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18356 word948 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18357 GND A9 word264 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18358 GND A4 word936 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18359 GND A4 word877 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18360 GND A8 word724 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18361 a_2162_n9004# a_2112_n66# a_1898_n9004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18362 GND A8 word163 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18363 a_2162_n85258# a_2112_n66# a_1898_n85258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18364 a_1238_n128142# A5 a_974_n128142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18365 word55 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18366 a_1766_n71626# A3 a_1370_n71626# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18367 GND A8 word104 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18368 a_1766_n80004# A3 a_1370_n80004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18369 a_1238_n119764# A5 a_842_n119764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18370 a_710_n89376# A7 a_446_n89376# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18371 a_446_n107978# A8 a_50_n107978# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18372 a_1766_n10282# A3 a_1502_n10282# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18373 GND A1 word156 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18374 word886 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18375 GND A1 word97 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18376 GND A6 word33 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18377 GND A2 word224 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18378 GND A7 word790 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18379 word971 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18380 GND A8 word651 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18381 word827 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18382 word491 a_2376_n66# a_2162_n69922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18383 GND A7 word346 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18384 GND A0 word756 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18385 a_50_n118912# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18386 a_446_n75034# A8 a_50_n75034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18387 a_1766_n57142# A3 a_1370_n57142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18388 GND A8 word721 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18389 a_1766_n48764# A3 a_1370_n48764# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18390 a_2294_n113374# A1 a_1898_n113374# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18391 a_1502_n128710# A4 a_1238_n128710# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18392 GND A7 word21 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18393 a_2294_n83270# A1 a_2030_n83270# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18394 GND A6 word186 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18395 a_1238_n110676# A5 a_974_n110676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18396 word782 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18397 a_710_n80288# A7 a_446_n80288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18398 GND A4 word711 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18399 word799 a_2376_n66# a_2162_n113658# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18400 word280 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18401 a_1370_n61828# a_1320_n66# a_1106_n61828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18402 word995 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18403 word860 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18404 GND A1 word205 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18405 word427 a_2376_n66# a_2162_n60834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18406 GND A7 word282 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18407 a_1502_n136662# A4 a_1238_n136662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18408 a_710_n124876# A7 a_314_n124876# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18409 a_974_n2046# A6 a_710_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18410 a_1370_n38966# a_1320_n66# a_1238_n38966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18411 word650 A0 a_2162_n92500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18412 GND A7 word612 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18413 GND A0 word1022 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18414 GND A8 word209 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18415 GND A7 word553 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18416 a_1766_n86536# A3 a_1502_n86536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18417 GND A1 word693 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18418 word117 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18419 GND A7 word121 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18420 a_2294_n142768# A1 a_1898_n142768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18421 word857 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18422 a_1766_n25192# A3 a_1370_n25192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18423 GND A1 word261 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18424 GND A7 word895 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18425 a_1502_n105138# A4 a_1106_n105138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18426 word989 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18427 word957 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18428 word605 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18429 word17 a_2376_n66# a_2294_n2614# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18430 GND A5 word16 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18431 a_842_n30304# a_792_n66# a_578_n30304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18432 a_974_n37404# A6 a_710_n37404# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18433 word887 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18434 GND A8 word145 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18435 word828 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18436 GND A1 word900 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18437 a_1370_n85116# a_1320_n66# a_1238_n85116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18438 a_50_n89802# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18439 a_1370_n76738# a_1320_n66# a_1238_n76738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18440 GND A8 word534 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18441 a_314_n40812# a_264_n66# a_182_n40812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18442 word591 a_2376_n66# a_2162_n84122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18443 word602 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18444 a_1370_n134248# a_1320_n66# a_1106_n134248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18445 a_50_n133112# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18446 GND A0 word738 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18447 a_1370_n125870# a_1320_n66# a_1106_n125870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18448 a_446_n1336# A8 a_182_n1336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18449 a_50_n124734# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18450 GND A7 word328 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18451 a_974_n8578# A6 a_710_n8578# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18452 GND A1 word468 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18453 a_1106_n35558# a_1056_n66# a_842_n35558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18454 a_578_n27606# a_528_n66# a_446_n27606# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18455 word1021 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18456 GND A5 word65 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18457 a_50_n80714# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18458 word380 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18459 GND A5 word768 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18460 word21 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18461 word5 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18462 GND A2 word592 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18463 GND A5 word926 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18464 a_578_n96902# a_528_n66# a_446_n96902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18465 a_1502_n142484# A4 a_1106_n142484# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18466 a_1370_n44788# a_1320_n66# a_1106_n44788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18467 a_1370_n53166# a_1320_n66# a_1106_n53166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18468 GND A0 word1004 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18469 GND A8 word250 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18470 GND A7 word594 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18471 a_1766_n7726# A3 a_1370_n7726# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18472 a_50_n101162# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18473 word158 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18474 word217 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18475 word307 a_2376_n66# a_2162_n43794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18476 a_182_n17808# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18477 a_314_n55722# a_264_n66# a_182_n55722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18478 word956 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18479 word914 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18480 GND A0 word902 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18481 GND A5 word704 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18482 GND A6 word434 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18483 a_446_n7868# A8 a_182_n7868# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18484 a_50_n139644# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18485 a_2030_n6022# A2 a_1634_n6022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18486 word43 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18487 a_446_n87388# A8 a_50_n87388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18488 GND A5 word975 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18489 word481 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18490 word212 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18491 a_974_n43226# A6 a_710_n43226# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18492 GND A1 word1000 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18493 GND A3 word945 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18494 word85 a_2376_n66# a_2294_n12270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18495 GND A6 word273 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18496 a_1106_n81282# a_1056_n66# a_974_n81282# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18497 word869 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18498 a_578_n64952# a_528_n66# a_314_n64952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18499 word945 a_2376_n66# a_2294_n134390# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18500 a_710_n6164# A7 a_446_n6164# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18501 a_50_n95624# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18502 word415 a_2376_n66# a_2162_n59130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18503 a_1370_n140070# a_1320_n66# a_1238_n140070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18504 word850 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18505 word774 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18506 a_842_n13264# a_792_n66# a_710_n13264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18507 a_50_n108120# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18508 a_1634_n8436# a_1584_n66# a_1370_n8436# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18509 a_2294_n9856# A1 a_1898_n9856# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18510 GND A0 word334 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18511 word573 a_2376_n66# a_2294_n81566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18512 GND A2 word697 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18513 word715 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18514 GND A2 word896 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18515 a_50_n130556# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18516 GND A7 word369 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18517 GND A1 word509 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18518 GND A4 word327 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18519 GND A4 word386 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18520 a_1370_n68076# a_1320_n66# a_1238_n68076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18521 word546 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18522 a_1106_n41380# a_1056_n66# a_974_n41380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18523 a_578_n33428# a_528_n66# a_446_n33428# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18524 a_1898_n15536# a_1848_n66# a_1634_n15536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18525 word471 a_2376_n66# a_2162_n67082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18526 a_1766_n98890# A3 a_1370_n98890# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18527 a_50_n107694# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18528 a_50_n116072# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18529 word10 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18530 a_182_n63532# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18531 GND A3 word167 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18532 a_314_n125302# a_264_n66# a_50_n125302# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18533 a_1106_n88240# a_1056_n66# a_842_n88240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18534 word716 A0 a_2294_n101872# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18535 a_314_n116924# a_264_n66# a_50_n116924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18536 GND A6 word539 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18537 word256 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18538 GND A2 word633 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18539 a_1502_n5312# A4 a_1106_n5312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18540 GND A4 word105 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18541 a_1898_n84832# a_1848_n66# a_1766_n84832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18542 a_842_n51036# a_792_n66# a_710_n51036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18543 a_974_n58136# A6 a_578_n58136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18544 word317 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18545 GND A7 word635 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18546 GND A0 word168 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18547 a_974_n80572# A6 a_710_n80572# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18548 a_1106_n96192# a_1056_n66# a_974_n96192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18549 a_182_n5454# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18550 a_182_n32008# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18551 a_314_n39108# a_264_n66# a_182_n39108# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18552 a_1502_n14116# A4 a_1106_n14116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18553 a_182_n23630# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18554 a_314_n61544# a_264_n66# a_182_n61544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18555 GND A4 word161 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18556 a_842_n89518# a_792_n66# a_710_n89518# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18557 word1014 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18558 word997 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18559 GND A4 word102 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18560 word879 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18561 a_842_n28174# a_792_n66# a_578_n28174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18562 a_1898_n53308# a_1848_n66# a_1766_n53308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18563 word529 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18564 word732 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18565 a_842_n142910# a_792_n66# a_578_n142910# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18566 word824 A0 a_2294_n117208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18567 a_50_n145466# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18568 word470 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18569 GND A0 word656 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18570 a_1502_n83412# A4 a_1238_n83412# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18571 word463 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18572 a_182_n31582# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18573 a_314_n38682# a_264_n66# a_182_n38682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18574 a_974_n40670# A6 a_710_n40670# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18575 a_50_n79010# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18576 GND A6 word314 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18577 a_578_n70774# a_528_n66# a_314_n70774# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18578 GND A3 word272 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18579 word524 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18580 a_1634_n5880# a_1584_n66# a_1502_n5880# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18581 word92 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18582 a_974_n26186# A6 a_578_n26186# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18583 a_1898_n99742# a_1848_n66# a_1634_n99742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18584 GND A2 word937 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18585 word587 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18586 word806 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18587 a_50_n78584# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18588 a_974_n95482# A6 a_578_n95482# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18589 a_1898_n21358# a_1848_n66# a_1766_n21358# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18590 a_182_n38540# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18591 a_1898_n4176# a_1848_n66# a_1634_n4176# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18592 a_1502_n29026# A4 a_1238_n29026# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18593 word304 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18594 word245 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18595 a_1502_n51462# A4 a_1106_n51462# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18596 a_314_n131124# a_264_n66# a_50_n131124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18597 a_1106_n134532# a_1056_n66# a_974_n134532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18598 a_1634_n126722# a_1584_n66# a_1370_n126722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18599 a_182_n60976# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18600 GND A4 word207 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18601 word262 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18602 a_1898_n68218# a_1848_n66# a_1634_n68218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18603 a_314_n122746# a_264_n66# a_50_n122746# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18604 word641 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18605 word297 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18606 a_1898_n59840# a_1848_n66# a_1766_n59840# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18607 word837 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18608 a_1898_n90654# a_1848_n66# a_1634_n90654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18609 GND A0 word702 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18610 GND A5 word146 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18611 word358 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18612 a_182_n46492# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18613 a_974_n55580# A6 a_578_n55580# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18614 GND A6 word419 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18615 a_578_n94062# a_528_n66# a_446_n94062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18616 word421 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18617 word880 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18618 GND A0 word150 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18619 a_1898_n67792# a_1848_n66# a_1634_n67792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18620 a_1238_n75602# A5 a_974_n75602# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18621 a_182_n2898# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18622 word629 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18623 word197 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18624 GND A0 word480 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18625 word570 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18626 word911 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18627 GND A0 word638 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18628 word692 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18629 word39 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18630 word504 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18631 word199 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18632 a_1370_n3466# a_1320_n66# a_1238_n3466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18633 a_1898_n36268# a_1848_n66# a_1634_n36268# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18634 a_842_n125870# a_792_n66# a_710_n125870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18635 word350 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18636 GND A3 word372 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18637 word409 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18638 word565 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18639 word98 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18640 a_314_n137656# a_264_n66# a_50_n137656# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18641 a_974_n100026# A6 a_578_n100026# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18642 a_1766_n103434# A3 a_1370_n103434# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18643 GND A6 word685 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18644 word687 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18645 word402 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18646 a_710_n40102# A7 a_314_n40102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18647 word179 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18648 GND A0 word26 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18649 a_1634_n13548# a_1584_n66# a_1370_n13548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18650 a_2030_n13832# A2 a_1766_n13832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18651 word847 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18652 word712 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18653 word569 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18654 word586 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18655 a_2162_n13122# a_2112_n66# a_2030_n13122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18656 word404 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18657 word667 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18658 a_2162_n136804# a_2112_n66# a_2030_n136804# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18659 GND A4 word680 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18660 word308 A0 a_2294_n43936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18661 word465 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18662 word303 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18663 a_1106_n131976# a_1056_n66# a_974_n131976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18664 a_1238_n4176# A5 a_974_n4176# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18665 word296 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18666 GND A3 word579 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18667 a_842_n102298# a_792_n66# a_578_n102298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18668 GND A6 word917 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18669 a_1238_n12128# A5 a_842_n12128# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18670 word237 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18671 a_1502_n95766# A4 a_1106_n95766# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18672 a_1766_n141206# A3 a_1502_n141206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18673 GND A3 word147 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18674 word206 A0 a_2162_n29452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18675 a_1766_n132828# A3 a_1502_n132828# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18676 a_2294_n11134# A1 a_1898_n11134# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18677 a_578_n69070# a_528_n66# a_314_n69070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18678 a_1634_n51320# a_1584_n66# a_1502_n51320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18679 a_2030_n51604# A2 a_1634_n51604# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18680 a_314_n114084# a_264_n66# a_50_n114084# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18681 a_2030_n111954# A2 a_1766_n111954# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18682 a_1106_n117492# a_1056_n66# a_974_n117492# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18683 GND A5 word517 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18684 GND A3 word418 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18685 a_2294_n49616# A1 a_1898_n49616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18686 word203 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18687 word670 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18688 a_1766_n118344# A3 a_1502_n118344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18689 a_2162_n42516# a_2112_n66# a_2030_n42516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18690 GND A3 word576 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18691 a_1766_n109966# A3 a_1502_n109966# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18692 a_2030_n28742# A2 a_1634_n28742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18693 a_710_n46634# A7 a_314_n46634# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18694 GND A8 word31 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18695 word361 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18696 word952 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18697 word501 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18698 word574 A0 a_2162_n81708# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18699 a_1238_n58562# A5 a_974_n58562# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18700 word510 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18701 GND A4 word514 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18702 word758 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18703 a_1898_n127006# a_1848_n66# a_1634_n127006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18704 word142 A0 a_2162_n20364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18705 word632 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18706 word78 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18707 word240 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18708 word562 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18709 a_842_n140070# a_792_n66# a_578_n140070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18710 a_446_n23914# A8 a_182_n23914# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18711 a_1898_n42090# a_1848_n66# a_1766_n42090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18712 word503 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18713 a_1634_n97754# a_1584_n66# a_1502_n97754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18714 GND A1 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18715 word472 A0 a_2294_n67224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18716 GND A3 word354 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18717 GND A9 word229 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18718 word881 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18719 a_710_n15110# A7 a_446_n15110# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18720 word80 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18721 a_2294_n40528# A1 a_1898_n40528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18722 a_314_n143478# a_264_n66# a_50_n143478# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18723 a_1766_n100878# A3 a_1502_n100878# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18724 GND A5 word134 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18725 word566 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18726 GND A5 word351 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18727 GND A3 word625 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18728 a_1238_n18660# A5 a_974_n18660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18729 GND A9 word127 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18730 word445 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18731 a_2030_n66514# A2 a_1766_n66514# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18732 a_710_n84406# A7 a_446_n84406# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18733 a_2162_n142626# a_2112_n66# a_2030_n142626# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18734 a_710_n14684# A7 a_446_n14684# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18735 word936 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18736 a_2162_n57426# a_2112_n66# a_2030_n57426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18737 word17 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18738 GND A5 word70 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18739 word120 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18740 word466 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18741 a_1634_n74182# a_1584_n66# a_1502_n74182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18742 word547 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18743 word615 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18744 GND A4 word619 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18745 a_2162_n119764# a_2112_n66# a_2030_n119764# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18746 word188 A0 a_2294_n26896# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18747 word183 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18748 word608 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18749 word176 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18750 GND A9 word393 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18751 GND A9 word334 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18752 a_2294_n55438# A1 a_1898_n55438# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18753 GND A3 word400 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18754 GND A1 word717 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18755 GND A6 word797 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18756 a_2030_n95908# A2 a_1766_n95908# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18757 word671 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18758 a_974_n112380# A6 a_710_n112380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18759 a_2030_n34564# A2 a_1766_n34564# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18760 a_710_n52456# A7 a_314_n52456# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18761 word325 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18762 GND A5 word397 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18763 word858 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18764 word301 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18765 a_1238_n64384# A5 a_842_n64384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18766 GND A8 word174 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18767 a_2162_n86820# a_2112_n66# a_2030_n86820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18768 word711 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18769 a_1238_n129704# A5 a_974_n129704# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18770 a_2162_n110676# a_2112_n66# a_2030_n110676# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18771 GND A7 word86 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18772 word550 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18773 a_2162_n25476# a_2112_n66# a_2030_n25476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18774 a_1766_n11844# A3 a_1370_n11844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18775 GND A7 word860 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18776 word454 A0 a_2162_n64668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18777 word982 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18778 word863 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18779 word390 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18780 a_2162_n94772# a_2112_n66# a_2030_n94772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18781 a_1634_n144898# a_1584_n66# a_1370_n144898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18782 a_2294_n114936# A1 a_2030_n114936# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18783 a_446_n15252# A8 a_182_n15252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18784 word79 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18785 word383 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18786 GND A7 word32 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18787 word793 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18788 GND A9 word168 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18789 GND A1 word924 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18790 a_1238_n120616# A5 a_842_n120616# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18791 GND A2 word291 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18792 a_710_n90228# A7 a_446_n90228# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18793 word761 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18794 GND A7 word857 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18795 GND A9 word109 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18796 a_2030_n141064# A2 a_1766_n141064# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18797 GND A4 word781 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18798 a_578_n134532# a_528_n66# a_314_n134532# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18799 a_2294_n23488# A1 a_1898_n23488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18800 a_710_n81850# A7 a_446_n81850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18801 a_2030_n63958# A2 a_1766_n63958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18802 GND A5 word663 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18803 word16 A0 a_2294_n2472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18804 GND A5 word604 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18805 word760 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18806 a_1238_n93778# A5 a_974_n93778# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18807 GND A6 word902 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18808 word918 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18809 GND A7 word293 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18810 a_1766_n139076# A3 a_1370_n139076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18811 a_974_n3608# A6 a_710_n3608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18812 word76 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18813 a_2294_n92784# A1 a_1898_n92784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18814 word767 a_2376_n66# a_2162_n109114# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18815 a_1634_n49190# a_1584_n66# a_1370_n49190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18816 a_2030_n49474# A2 a_1634_n49474# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18817 word507 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18818 word647 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18819 GND A1 word921 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18820 a_1370_n48906# a_1320_n66# a_1238_n48906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18821 word731 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18822 word288 A0 a_2294_n41096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18823 a_578_n103008# a_528_n66# a_446_n103008# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18824 a_1898_n139360# a_1848_n66# a_1766_n139360# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18825 a_2162_n125586# a_2112_n66# a_2030_n125586# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18826 word757 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18827 word986 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18828 word927 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18829 a_1766_n35132# A3 a_1370_n35132# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18830 GND A1 word272 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18831 GND A3 word500 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18832 GND A9 word375 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18833 GND A9 word47 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18834 a_1106_n16104# a_1056_n66# a_842_n16104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18835 GND A2 word498 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18836 word703 a_2376_n66# a_2162_n100026# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18837 a_2294_n138224# A1 a_1898_n138224# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18838 a_2294_n129846# A1 a_2030_n129846# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18839 a_2030_n40386# A2 a_1634_n40386# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18840 a_578_n102582# a_528_n66# a_446_n102582# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18841 word766 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18842 GND A1 word56 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18843 word125 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18844 word184 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18845 word488 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18846 GND A8 word215 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18847 word898 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18848 a_1502_n114652# A4 a_1106_n114652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18849 a_2162_n31298# a_2112_n66# a_2030_n31298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18850 a_2294_n38398# A1 a_1898_n38398# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18851 a_2030_n78868# A2 a_1634_n78868# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18852 a_710_n111244# A7 a_314_n111244# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18853 a_1370_n16956# a_1320_n66# a_1106_n16956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18854 a_1370_n25334# a_1320_n66# a_1106_n25334# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18855 word1023 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18856 a_1370_n135810# a_1320_n66# a_1106_n135810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18857 GND A0 word808 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18858 GND A8 word113 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18859 a_446_n82418# A8 a_50_n82418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18860 a_1766_n64526# A3 a_1502_n64526# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18861 a_2162_n69780# a_2112_n66# a_2030_n69780# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18862 word111 a_2376_n66# a_2162_n15962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18863 a_2294_n120758# A1 a_2030_n120758# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18864 a_446_n12696# A8 a_182_n12696# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18865 a_446_n21074# A8 a_182_n21074# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18866 GND A6 word42 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18867 GND A2 word115 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18868 GND A8 word601 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18869 GND A9 word150 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18870 a_1370_n143762# a_1320_n66# a_1106_n143762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18871 a_578_n140354# a_528_n66# a_314_n140354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18872 a_578_n131976# a_528_n66# a_314_n131976# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18873 GND A5 word645 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18874 word695 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18875 a_2294_n342# A1 a_2030_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18876 a_446_n81992# A8 a_50_n81992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18877 GND A9 word480 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18878 GND A6 word136 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18879 GND A2 word603 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18880 GND A9 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18881 GND A1 word804 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18882 a_446_n100168# A8 a_50_n100168# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18883 a_1238_n103576# A5 a_842_n103576# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18884 GND A1 word745 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18885 GND A2 word171 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18886 a_710_n73188# A7 a_446_n73188# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18887 a_1370_n63106# a_1320_n66# a_1106_n63106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18888 word749 a_2376_n66# a_2294_n106558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18889 word506 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18890 word447 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18891 word810 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18892 a_1370_n112238# a_1320_n66# a_1238_n112238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18893 a_50_n111102# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18894 word377 a_2376_n66# a_2294_n53734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18895 a_1766_n93920# A3 a_1370_n93920# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18896 a_1370_n103860# a_1320_n66# a_1238_n103860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18897 a_1502_n129562# A4 a_1238_n129562# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18898 a_710_n126154# A7 a_314_n126154# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18899 a_50_n102724# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18900 GND A1 word313 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18901 GND A1 word372 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18902 a_710_n117776# A7 a_314_n117776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18903 GND A4 word131 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18904 a_1766_n32576# A3 a_1502_n32576# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18905 GND A8 word57 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18906 word984 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18907 GND A0 word972 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18908 GND A5 word774 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18909 GND A5 word715 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18910 word600 A0 a_2294_n85400# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18911 a_446_n97328# A8 a_50_n97328# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18912 word1009 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18913 a_446_n88950# A8 a_50_n88950# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18914 a_2294_n144046# A1 a_1898_n144046# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18915 word155 a_2376_n66# a_2162_n22210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18916 GND A3 word1015 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18917 word939 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18918 GND A0 word74 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18919 GND A2 word378 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18920 word1015 a_2376_n66# a_2162_n144330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18921 GND A4 word868 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18922 a_1502_n120474# A4 a_1238_n120474# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18923 a_710_n7726# A7 a_446_n7726# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18924 word555 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18925 a_2030_n84690# A2 a_1766_n84690# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18926 word920 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18927 a_1370_n22778# a_1320_n66# a_1238_n22778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18928 a_1370_n31156# a_1320_n66# a_1238_n31156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18929 word643 a_2376_n66# a_2162_n91506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18930 a_842_n14826# a_792_n66# a_710_n14826# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18931 GND A8 word95 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18932 GND A8 word154 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18933 word837 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18934 GND A1 word909 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18935 a_1238_n118486# A5 a_842_n118486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18936 word211 a_2376_n66# a_2162_n30162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18937 a_1106_n59982# a_1056_n66# a_974_n59982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18938 a_446_n106700# A8 a_50_n106700# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18939 a_1766_n61970# A3 a_1370_n61970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18940 a_710_n88098# A7 a_446_n88098# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18941 GND A1 word88 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18942 word552 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18943 word801 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18944 word818 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18945 a_1106_n51320# a_1056_n66# a_842_n51320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18946 word541 a_2376_n66# a_2294_n77022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18947 GND A8 word642 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18948 a_1370_n127148# a_1320_n66# a_1106_n127148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18949 word759 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18950 a_50_n126012# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18951 GND A7 word278 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18952 GND A7 word337 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18953 GND A8 word583 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18954 a_50_n117634# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18955 a_2294_n112096# A1 a_1898_n112096# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18956 word786 A0 a_2162_n111812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18957 a_974_n21216# A6 a_578_n21216# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18958 GND A1 word576 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18959 a_2030_n626# A2 a_1766_n626# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18960 GND A6 word177 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18961 GND A1 word845 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18962 GND A3 word790 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18963 a_1106_n50894# a_1056_n66# a_842_n50894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18964 word971 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18965 word330 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18966 a_50_n73614# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18967 a_1106_n97754# a_1056_n66# a_974_n97754# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18968 GND A2 word483 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18969 GND A4 word973 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18970 a_710_n123598# A7 a_314_n123598# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18971 GND A4 word172 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18972 GND A4 word231 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18973 GND A7 word544 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18974 GND A0 word954 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18975 a_842_n29736# a_792_n66# a_578_n29736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18976 GND A8 word200 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18977 GND A1 word684 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18978 word743 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18979 word257 a_2376_n66# a_2294_n36694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18980 a_1766_n85258# A3 a_1370_n85258# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18981 GND A1 word625 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18982 a_182_n41522# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18983 a_314_n48622# a_264_n66# a_182_n48622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18984 GND A6 word384 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18985 GND A6 word443 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18986 GND A8 word688 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18987 a_446_n9146# A8 a_182_n9146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18988 word946 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18989 word596 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18990 GND A5 word7 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18991 word103 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X18992 word819 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18993 a_2162_n5170# a_2112_n66# a_2030_n5170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18994 word895 a_2376_n66# a_2162_n127290# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18995 a_1238_n484# A5 a_974_n484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18996 a_578_n57852# a_528_n66# a_314_n57852# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18997 a_1370_n75460# a_1320_n66# a_1238_n75460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X18998 a_50_n88524# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X18999 a_842_n67508# a_792_n66# a_578_n67508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19000 word859 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19001 GND A4 word11 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19002 GND A5 word2 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19003 word523 a_2376_n66# a_2162_n74466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19004 GND A0 word788 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19005 a_1898_n5738# a_1848_n66# a_1766_n5738# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19006 word374 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19007 GND A7 word319 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19008 a_974_n7300# A6 a_710_n7300# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19009 a_50_n123456# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19010 word315 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19011 a_1502_n61402# A4 a_1106_n61402# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19012 GND A0 word442 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19013 a_182_n70916# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19014 GND A1 word400 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19015 word367 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19016 word308 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19017 a_1106_n34280# a_1056_n66# a_842_n34280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19018 a_842_n106416# a_792_n66# a_578_n106416# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19019 a_578_n26328# a_528_n66# a_446_n26328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19020 GND A6 word159 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19021 a_182_n56432# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19022 GND A3 word117 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19023 word371 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19024 a_314_n118202# a_264_n66# a_50_n118202# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19025 GND A6 word548 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19026 a_2294_n2046# A1 a_1898_n2046# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19027 a_314_n109824# a_264_n66# a_50_n109824# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19028 word491 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19029 GND A0 word220 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19030 a_578_n95624# a_528_n66# a_446_n95624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19031 GND A2 word723 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19032 word701 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19033 GND A7 word585 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19034 a_842_n35558# a_792_n66# a_578_n35558# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19035 a_974_n73472# A6 a_710_n73472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19036 a_1106_n89092# a_1056_n66# a_842_n89092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19037 word981 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19038 a_1766_n91080# A3 a_1502_n91080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19039 word1006 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19040 a_182_n16530# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19041 word90 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19042 word149 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19043 GND A4 word484 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19044 word947 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19045 a_314_n54444# a_264_n66# a_182_n54444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19046 a_1898_n46208# a_1848_n66# a_1766_n46208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19047 GND A6 word425 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19048 word427 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19049 word770 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19050 a_50_n138366# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19051 word34 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19052 word479 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19053 GND A0 word606 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19054 word987 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19055 a_446_n6590# A8 a_182_n6590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19056 a_50_n129988# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19057 word637 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19058 word932 A0 a_2294_n132544# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19059 word472 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19060 a_182_n24482# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19061 word413 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19062 word917 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19063 a_578_n72052# a_528_n66# a_314_n72052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19064 GND A6 word264 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19065 word639 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19066 word826 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19067 a_50_n94346# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19068 a_578_n63674# a_528_n66# a_314_n63674# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19069 a_842_n143762# a_792_n66# a_578_n143762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19070 a_50_n85968# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19071 GND A3 word21 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19072 word476 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19073 a_974_n19086# A6 a_578_n19086# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19074 word710 A0 a_2162_n101020# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19075 word756 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19076 a_50_n120900# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19077 GND A1 word500 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19078 word537 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19079 a_1106_n141916# a_1056_n66# a_842_n141916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19080 word11 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19081 GND A4 word259 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19082 a_578_n32150# a_528_n66# a_446_n32150# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19083 word254 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19084 a_1634_n69922# a_1584_n66# a_1502_n69922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19085 a_842_n103860# a_792_n66# a_578_n103860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19086 a_314_n69354# a_264_n66# a_182_n69354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19087 a_182_n53876# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19088 a_182_n62254# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19089 a_314_n115646# a_264_n66# a_50_n115646# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19090 a_314_n124024# a_264_n66# a_50_n124024# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19091 a_1634_n119622# a_1584_n66# a_1502_n119622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19092 GND A6 word530 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19093 GND A3 word646 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19094 a_182_n39392# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19095 a_1238_n21642# A5 a_974_n21642# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19096 word963 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19097 word1022 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19098 GND A0 word100 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19099 a_1634_n60834# a_1584_n66# a_1502_n60834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19100 GND A4 word584 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19101 word830 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19102 a_182_n4176# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19103 word212 A0 a_2294_n30304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19104 GND A4 word525 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19105 a_314_n51888# a_264_n66# a_182_n51888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19106 a_314_n60266# a_264_n66# a_182_n60266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19107 a_842_n88240# a_792_n66# a_710_n88240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19108 a_1634_n110534# a_1584_n66# a_1502_n110534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19109 a_1898_n52030# a_1848_n66# a_1634_n52030# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19110 word669 a_2376_n66# a_2294_n95198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19111 a_50_n144188# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19112 a_1634_n37972# a_1584_n66# a_1502_n37972# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19113 a_1502_n82134# A4 a_1238_n82134# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19114 GND A0 word588 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19115 a_1502_n73756# A4 a_1238_n73756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19116 word454 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19117 a_1898_n29168# a_1848_n66# a_1634_n29168# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19118 a_842_n127148# a_792_n66# a_710_n127148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19119 a_842_n118770# a_792_n66# a_710_n118770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19120 GND A3 word263 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19121 a_182_n68786# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19122 a_50_n91790# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19123 a_2294_n27606# A1 a_2030_n27606# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19124 a_1502_n59272# A4 a_1106_n59272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19125 word696 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19126 a_2030_n136804# A2 a_1766_n136804# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19127 a_2162_n20506# a_2112_n66# a_1898_n20506# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19128 word129 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19129 a_1898_n98464# a_1848_n66# a_1766_n98464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19130 word797 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19131 GND A5 word201 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19132 word287 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19133 word578 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19134 word738 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19135 a_1238_n36552# A5 a_974_n36552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19136 GND A4 word300 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19137 word355 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19138 GND A4 word359 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19139 word519 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19140 word477 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19141 a_2294_n96902# A1 a_2030_n96902# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19142 a_1634_n84122# a_1584_n66# a_1502_n84122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19143 word617 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19144 a_1898_n20080# a_1848_n66# a_1634_n20080# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19145 a_1502_n19370# A4 a_1238_n19370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19146 word258 A0 a_2162_n36836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19147 GND A9 word74 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19148 a_314_n66798# a_264_n66# a_182_n66798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19149 a_1502_n50184# A4 a_1106_n50184# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19150 a_314_n121468# a_264_n66# a_50_n121468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19151 word415 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19152 a_1106_n133254# a_1056_n66# a_974_n133254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19153 a_1106_n124876# a_1056_n66# a_842_n124876# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19154 word194 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19155 word288 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19156 word246 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19157 GND A3 word529 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19158 a_1502_n1478# A4 a_1238_n1478# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19159 word187 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19160 GND A3 word470 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19161 a_1502_n88666# A4 a_1106_n88666# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19162 a_1502_n97044# A4 a_1106_n97044# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19163 GND A6 word808 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19164 word255 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19165 a_1766_n125728# A3 a_1370_n125728# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19166 a_2030_n44504# A2 a_1634_n44504# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19167 GND A5 word467 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19168 a_2030_n104854# A2 a_1766_n104854# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19169 word471 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19170 word1004 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19171 a_1238_n74324# A5 a_974_n74324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19172 a_1238_n65946# A5 a_842_n65946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19173 word620 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19174 word722 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19175 a_2294_n64952# A1 a_2030_n64952# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19176 a_974_n130272# A6 a_578_n130272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19177 a_710_n39534# A7 a_314_n39534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19178 word252 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19179 word451 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19180 word524 A0 a_2294_n74608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19181 word902 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19182 GND A9 word12 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19183 a_1634_n52172# a_1584_n66# a_1502_n52172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19184 a_2162_n106132# a_2112_n66# a_2030_n106132# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19185 word683 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19186 word767 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19187 GND A0 word20 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19188 word30 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19189 word92 A0 a_2294_n13264# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19190 word190 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19191 word495 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19192 a_1898_n133964# a_1848_n66# a_1634_n133964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19193 word676 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19194 a_1634_n99032# a_1584_n66# a_1370_n99032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19195 a_446_n16814# A8 a_182_n16814# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19196 GND A3 word304 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19197 a_1502_n65094# A4 a_1238_n65094# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19198 GND A9 word179 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19199 word831 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19200 GND A3 word245 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19201 a_314_n136378# a_264_n66# a_50_n136378# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19202 a_2030_n142626# A2 a_1634_n142626# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19203 a_314_n128000# a_264_n66# a_50_n128000# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19204 word678 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19205 GND A6 word913 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19206 a_2162_n64810# a_2112_n66# a_1898_n64810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19207 a_1106_n6732# a_1056_n66# a_974_n6732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19208 a_710_n77306# A7 a_446_n77306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19209 a_1634_n59130# a_1584_n66# a_1370_n59130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19210 a_2030_n59414# A2 a_1766_n59414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19211 word577 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19212 a_2030_n119764# A2 a_1634_n119764# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19213 a_1634_n81566# a_1584_n66# a_1370_n81566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19214 word974 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19215 GND A2 word35 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19216 word358 A0 a_2162_n51036# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19217 a_1634_n131266# a_1584_n66# a_1370_n131266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19218 word235 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19219 a_2162_n72762# a_2112_n66# a_1898_n72762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19220 a_2294_n79862# A1 a_2030_n79862# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19221 a_2294_n101304# A1 a_2030_n101304# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19222 word228 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19223 word138 A0 a_2162_n19796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19224 a_2030_n50326# A2 a_1766_n50326# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19225 word558 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19226 a_2030_n110676# A2 a_1634_n110676# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19227 GND A5 word449 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19228 word126 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19229 a_2030_n88808# A2 a_1766_n88808# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19230 a_710_n112806# A7 a_314_n112806# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19231 GND A9 word501 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19232 GND A9 word442 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19233 a_1766_n117066# A3 a_1370_n117066# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19234 a_2162_n32860# a_2112_n66# a_1898_n32860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19235 word275 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19236 a_2294_n39960# A1 a_2030_n39960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19237 a_2294_n70774# A1 a_2030_n70774# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19238 GND A8 word22 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19239 word352 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19240 a_710_n36978# A7 a_314_n36978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19241 a_710_n45356# A7 a_314_n45356# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19242 a_1634_n27180# a_1584_n66# a_1370_n27180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19243 a_2030_n27464# A2 a_1766_n27464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19244 GND A5 word347 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19245 word433 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19246 GND A8 word124 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19247 word749 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19248 word251 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19249 a_1238_n57284# A5 a_974_n57284# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19250 word181 a_2376_n66# a_2294_n25902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19251 word623 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19252 a_446_n22636# A8 a_182_n22636# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19253 a_446_n31014# A8 a_182_n31014# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19254 GND A1 word117 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19255 word494 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19256 GND A6 word53 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19257 word435 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19258 GND A7 word810 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19259 word404 A0 a_2294_n57568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19260 GND A9 word220 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19261 a_314_n142200# a_264_n66# a_50_n142200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19262 GND A8 word741 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19263 a_1634_n137798# a_1584_n66# a_1502_n137798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19264 word813 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19265 a_578_n141916# a_528_n66# a_314_n141916# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19266 a_2294_n116214# A1 a_2030_n116214# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19267 a_446_n91932# A8 a_50_n91932# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19268 GND A3 word675 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19269 GND A7 word41 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19270 GND A5 word283 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19271 a_2294_n86110# A1 a_1898_n86110# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19272 GND A6 word954 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19273 GND A7 word807 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19274 GND A7 word866 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19275 a_1238_n113516# A5 a_974_n113516# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19276 GND A2 word241 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19277 a_2030_n65236# A2 a_1634_n65236# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19278 a_710_n83128# A7 a_446_n83128# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19279 a_446_n101730# A8 a_50_n101730# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19280 a_2030_n125586# A2 a_1766_n125586# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19281 a_578_n127432# a_528_n66# a_314_n127432# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19282 a_710_n74750# A7 a_446_n74750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19283 word1015 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19284 a_1238_n95056# A5 a_974_n95056# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19285 a_2162_n141348# a_2112_n66# a_2030_n141348# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19286 a_2162_n132970# a_2112_n66# a_1898_n132970# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19287 GND A0 word712 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19288 a_2162_n47770# a_2112_n66# a_1898_n47770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19289 a_2162_n56148# a_2112_n66# a_2030_n56148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19290 a_2294_n94062# A1 a_1898_n94062# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19291 word457 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19292 GND A8 word68 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19293 word670 A0 a_2162_n95340# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19294 word936 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19295 word877 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19296 a_1370_n121752# a_1320_n66# a_1238_n121752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19297 a_1766_n28032# A3 a_1502_n28032# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19298 GND A9 word56 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19299 GND A3 word450 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19300 GND A9 word325 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19301 GND A6 word788 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19302 a_2294_n54160# A1 a_1898_n54160# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19303 GND A2 word448 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19304 a_2030_n94630# A2 a_1634_n94630# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19305 GND A0 a_2376_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X19306 a_710_n42800# A7 a_314_n42800# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19307 a_2030_n33286# A2 a_1634_n33286# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19308 a_710_n51178# A7 a_314_n51178# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19309 word351 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19310 GND A5 word388 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19311 GND A8 word165 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19312 GND A8 word224 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19313 word281 a_2376_n66# a_2294_n40102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19314 GND A2 word346 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19315 a_1106_n69922# a_1056_n66# a_842_n69922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19316 a_1238_n128426# A5 a_974_n128426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19317 GND A7 word77 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19318 a_710_n89660# A7 a_446_n89660# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19319 GND A1 word217 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19320 a_1370_n18234# a_1320_n66# a_1106_n18234# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19321 word622 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19322 word973 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19323 word829 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19324 GND A7 word348 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19325 GND A0 word758 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19326 word914 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19327 GND A8 word653 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19328 a_446_n75318# A8 a_50_n75318# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19329 a_1766_n57426# A3 a_1370_n57426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19330 GND A8 word221 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19331 GND A8 word723 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19332 GND A1 word976 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19333 GND A7 word23 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19334 a_1238_n110960# A5 a_974_n110960# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19335 word784 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19336 GND A8 word551 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19337 GND A9 word100 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19338 GND A2 word282 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19339 a_1106_n60834# a_1056_n66# a_974_n60834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19340 a_2030_n71058# A2 a_1766_n71058# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19341 GND A4 word713 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19342 a_578_n133254# a_528_n66# a_314_n133254# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19343 a_2030_n62680# A2 a_1634_n62680# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19344 GND A5 word595 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19345 GND A5 word654 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19346 a_446_n74892# A8 a_50_n74892# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19347 a_2294_n69070# A1 a_1898_n69070# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19348 GND A2 word553 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19349 a_1238_n92500# A5 a_974_n92500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19350 GND A7 word284 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19351 a_1502_n136946# A4 a_1238_n136946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19352 a_974_n2330# A6 a_710_n2330# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19353 GND A2 word121 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19354 GND A1 word424 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19355 GND A3 word916 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19356 a_2030_n48196# A2 a_1766_n48196# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19357 word397 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19358 word895 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19359 word857 a_2376_n66# a_2294_n121894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19360 word760 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19361 word327 a_2376_n66# a_2162_n46634# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19362 a_1766_n86820# A3 a_1502_n86820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19363 a_50_n104002# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19364 GND A7 word123 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19365 a_710_n119054# A7 a_314_n119054# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19366 a_1766_n25476# A3 a_1370_n25476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19367 GND A5 word724 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19368 a_446_n34990# A8 a_182_n34990# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19369 word550 A0 a_2162_n78300# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19370 GND A9 word38 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19371 word959 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19372 GND A7 word611 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19373 a_2294_n128568# A1 a_2030_n128568# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19374 a_578_n20932# a_528_n66# a_446_n20932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19375 word175 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19376 GND A5 word18 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19377 word105 a_2376_n66# a_2294_n15110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19378 GND A1 word1020 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19379 GND A3 word965 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19380 GND A7 word69 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19381 GND A2 word387 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19382 word889 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19383 word965 a_2376_n66# a_2294_n137230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19384 GND A5 word721 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19385 a_710_n9004# A7 a_446_n9004# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19386 GND A2 word328 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19387 a_2030_n77590# A2 a_1766_n77590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19388 a_578_n139786# a_528_n66# a_314_n139786# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19389 a_1502_n104996# A4 a_1106_n104996# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19390 word604 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19391 word1014 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19392 GND A0 word858 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19393 a_842_n16104# a_792_n66# a_710_n16104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19394 word593 a_2376_n66# a_2294_n84406# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19395 a_446_n1620# A8 a_182_n1620# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19396 a_446_n81140# A8 a_50_n81140# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19397 GND A0 word512 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19398 GND A1 word529 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19399 word161 a_2376_n66# a_2294_n23062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19400 a_1766_n54870# A3 a_1502_n54870# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19401 word1021 a_2376_n66# a_2294_n145182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19402 word751 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19403 a_1106_n44220# a_1056_n66# a_974_n44220# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19404 a_1370_n84974# a_1320_n66# a_1238_n84974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19405 a_1370_n93352# a_1320_n66# a_1238_n93352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19406 word1023 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19407 GND A8 word592 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19408 GND A8 word533 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19409 word926 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19410 a_1898_n40812# a_1848_n66# a_1634_n40812# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19411 word791 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19412 word441 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19413 word736 A0 a_2294_n104712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19414 a_578_n130698# a_528_n66# a_314_n130698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19415 word23 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19416 GND A5 word987 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19417 GND A5 word770 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19418 a_2294_n3608# A1 a_2030_n3608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19419 GND A2 word594 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19420 a_1106_n52172# a_1056_n66# a_842_n52172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19421 a_1238_n102298# A5 a_842_n102298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19422 GND A3 word740 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19423 a_1502_n142768# A4 a_1106_n142768# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19424 GND A2 word793 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19425 a_1106_n43794# a_1056_n66# a_974_n43794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19426 a_578_n35842# a_528_n66# a_446_n35842# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19427 a_1370_n53450# a_1320_n66# a_1106_n53450# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19428 a_1106_n99032# a_1056_n66# a_974_n99032# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19429 a_50_n101446# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19430 a_710_n116498# A7 a_314_n116498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19431 word1017 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19432 a_1502_n128284# A4 a_1238_n128284# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19433 a_1634_n1762# a_1584_n66# a_1502_n1762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19434 GND A1 word304 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19435 GND A1 word245 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19436 GND A0 word904 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19437 a_50_n139928# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19438 a_2030_n6306# A2 a_1634_n6306# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19439 a_446_n96050# A8 a_50_n96050# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19440 a_1766_n78158# A3 a_1502_n78158# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19441 word998 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19442 word207 a_2376_n66# a_2162_n29594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19443 a_2294_n134390# A1 a_2030_n134390# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19444 a_182_n34422# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19445 word216 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19446 a_974_n43510# A6 a_710_n43510# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19447 GND A6 word393 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19448 a_1370_n99884# a_1320_n66# a_1106_n99884# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19449 GND A8 word697 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19450 a_1238_n140070# A5 a_842_n140070# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19451 a_1106_n81566# a_1056_n66# a_974_n81566# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19452 word930 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19453 GND A2 word369 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19454 a_1898_n55722# a_1848_n66# a_1766_n55722# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19455 GND A4 word800 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19456 a_710_n6448# A7 a_446_n6448# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19457 a_50_n95908# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19458 GND A3 word32 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19459 a_842_n13548# a_792_n66# a_710_n13548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19460 a_1634_n8720# a_1584_n66# a_1370_n8720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19461 a_1370_n21500# a_1320_n66# a_1238_n21500# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19462 word575 a_2376_n66# a_2162_n81850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19463 GND A2 word699 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19464 GND A2 word898 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19465 a_50_n130840# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19466 word769 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19467 GND A4 word329 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19468 a_1370_n90796# a_1320_n66# a_1106_n90796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19469 a_974_n98322# A6 a_578_n98322# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19470 GND A8 word633 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19471 word473 a_2376_n66# a_2294_n67366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19472 a_842_n82844# a_792_n66# a_710_n82844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19473 a_50_n116356# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19474 a_1898_n15820# a_1848_n66# a_1634_n15820# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19475 GND A7 word269 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19476 a_182_n63816# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19477 a_50_n107978# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19478 GND A0 word392 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19479 GND A1 word409 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19480 a_1502_n45924# A4 a_1238_n45924# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19481 word317 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19482 a_1106_n27180# a_1056_n66# a_974_n27180# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19483 GND A2 word635 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19484 word258 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19485 a_578_n19228# a_528_n66# a_446_n19228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19486 GND A6 word168 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19487 word956 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19488 a_842_n121752# a_792_n66# a_710_n121752# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19489 a_182_n49332# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19490 a_1898_n23772# a_1848_n66# a_1766_n23772# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19491 a_974_n58420# A6 a_578_n58420# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19492 a_842_n51320# a_792_n66# a_710_n51320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19493 GND A0 word170 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19494 a_974_n80856# A6 a_710_n80856# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19495 a_1106_n96476# a_1056_n66# a_974_n96476# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19496 GND A6 word656 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19497 GND A4 word964 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19498 a_182_n5738# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19499 a_314_n70206# a_264_n66# a_182_n70206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19500 a_314_n61828# a_264_n66# a_182_n61828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19501 GND A4 word104 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19502 GND A4 word163 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19503 word63 a_2376_n66# a_2162_n9146# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19504 a_842_n28458# a_792_n66# a_578_n28458# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19505 GND A7 word535 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19506 a_974_n57994# A6 a_578_n57994# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19507 GND A0 word658 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19508 word734 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19509 a_2030_n3750# A2 a_1634_n3750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19510 a_842_n50894# a_792_n66# a_710_n50894# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19511 a_314_n47344# a_264_n66# a_182_n47344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19512 GND A0 word226 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19513 GND A4 word651 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19514 a_182_n31866# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19515 a_314_n38966# a_264_n66# a_182_n38966# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19516 a_182_n40244# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19517 a_1502_n13974# A4 a_1106_n13974# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19518 a_1106_n105422# a_1056_n66# a_842_n105422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19519 word436 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19520 GND A4 word66 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19521 GND A0 word556 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19522 word878 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19523 a_1502_n69212# A4 a_1106_n69212# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19524 word882 A0 a_2162_n125444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19525 a_182_n17382# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19526 GND A0 word46 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19527 word94 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19528 a_974_n26470# A6 a_578_n26470# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19529 word867 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19530 GND A2 word939 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19531 word808 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19532 word648 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19533 a_578_n56574# a_528_n66# a_314_n56574# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19534 a_1898_n38682# a_1848_n66# a_1634_n38682# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19535 GND A4 word429 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19536 word589 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19537 a_842_n136662# a_792_n66# a_578_n136662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19538 a_50_n87246# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19539 a_842_n66230# a_792_n66# a_578_n66230# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19540 a_50_n78868# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19541 word155 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19542 word582 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19543 a_974_n95766# A6 a_578_n95766# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19544 GND A6 word702 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19545 a_50_n122178# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19546 a_1898_n4460# a_1848_n66# a_1634_n4460# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19547 a_1502_n29310# A4 a_1238_n29310# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19548 GND A0 word492 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19549 a_50_n113800# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19550 a_1634_n15962# a_1584_n66# a_1502_n15962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19551 GND A4 word268 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19552 a_1502_n60124# A4 a_1106_n60124# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19553 a_1502_n51746# A4 a_1106_n51746# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19554 a_314_n131408# a_264_n66# a_50_n131408# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19555 word643 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19556 word358 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19557 a_1106_n134816# a_1056_n66# a_974_n134816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19558 GND A4 word426 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19559 word299 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19560 word839 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19561 a_578_n25050# a_528_n66# a_446_n25050# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19562 GND A6 word150 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19563 word421 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19564 word211 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19565 a_1898_n90938# a_1848_n66# a_1634_n90938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19566 a_842_n105138# a_792_n66# a_578_n105138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19567 word152 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19568 word997 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19569 a_182_n55154# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19570 a_1502_n37262# A4 a_1238_n37262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19571 a_182_n46776# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19572 a_1502_n28884# A4 a_1238_n28884# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19573 a_314_n130982# a_264_n66# a_50_n130982# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19574 word482 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19575 a_578_n94346# a_528_n66# a_446_n94346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19576 GND A2 word714 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19577 word692 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19578 word983 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19579 GND A3 word596 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19580 a_842_n34280# a_792_n66# a_578_n34280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19581 word199 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19582 word322 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19583 word381 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19584 word972 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19585 a_974_n131834# A6 a_578_n131834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19586 word775 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19587 a_1766_n5170# A3 a_1502_n5170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19588 word45 a_2376_n66# a_2294_n6590# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19589 word357 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19590 a_1634_n53734# a_1584_n66# a_1370_n53734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19591 word913 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19592 word694 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19593 a_314_n53166# a_264_n66# a_182_n53166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19594 word162 A0 a_2162_n23204# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19595 word938 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19596 a_314_n44788# a_264_n66# a_182_n44788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19597 word98 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19598 word687 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19599 a_1898_n143904# a_1848_n66# a_1766_n143904# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19600 word619 a_2376_n66# a_2162_n88098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19601 a_1370_n3750# a_1320_n66# a_1238_n3750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19602 a_50_n137088# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19603 GND A3 word374 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19604 GND A0 word538 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19605 word919 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19606 GND A1 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19607 a_1502_n75034# A4 a_1238_n75034# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19608 word569 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19609 word864 A0 a_2294_n122888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19610 word66 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19611 a_314_n137940# a_264_n66# a_50_n137940# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19612 word586 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19613 word404 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19614 a_1634_n22210# a_1584_n66# a_1370_n22210# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19615 a_842_n89092# a_792_n66# a_710_n89092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19616 word849 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19617 a_578_n62396# a_528_n66# a_314_n62396# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19618 a_842_n142484# a_792_n66# a_578_n142484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19619 a_50_n93068# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19620 GND A7 word836 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19621 a_2030_n129704# A2 a_1766_n129704# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19622 a_50_n84690# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19623 GND A3 word371 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19624 a_2294_n42942# A1 a_1898_n42942# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19625 a_710_n17524# A7 a_446_n17524# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19626 word97 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19627 word747 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19628 GND A2 word819 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19629 a_1634_n21784# a_1584_n66# a_1370_n21784# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19630 word237 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19631 word528 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19632 a_1238_n29452# A5 a_842_n29452# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19633 word486 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19634 a_842_n49190# a_792_n66# a_710_n49190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19635 a_1634_n77022# a_1584_n66# a_1370_n77022# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19636 a_1898_n120332# a_1848_n66# a_1634_n120332# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19637 a_1238_n4460# A5 a_974_n4460# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19638 word298 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19639 a_314_n68076# a_264_n66# a_182_n68076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19640 GND A3 word149 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19641 word208 A0 a_2294_n29736# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19642 a_1502_n43084# A4 a_1106_n43084# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19643 a_1106_n126154# a_1056_n66# a_842_n126154# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19644 a_182_n52598# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19645 a_314_n59698# a_264_n66# a_182_n59698# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19646 word203 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19647 a_314_n114368# a_264_n66# a_50_n114368# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19648 a_2030_n120616# A2 a_1766_n120616# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19649 a_1106_n117776# a_1056_n66# a_974_n117776# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19650 a_1898_n73898# a_1848_n66# a_1766_n73898# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19651 a_578_n91790# a_528_n66# a_446_n91790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19652 GND A6 word817 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19653 GND A5 word87 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19654 GND A3 word420 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19655 a_1238_n20364# A5 a_974_n20364# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19656 word205 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19657 word691 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19658 a_2030_n106132# A2 a_1634_n106132# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19659 a_1766_n118628# A3 a_1502_n118628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19660 a_974_n115220# A6 a_710_n115220# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19661 a_1238_n11986# A5 a_842_n11986# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19662 word363 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19663 word1013 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19664 a_710_n46918# A7 a_314_n46918# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19665 word503 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19666 word954 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19667 a_2294_n10992# A1 a_1898_n10992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19668 a_1238_n67224# A5 a_842_n67224# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19669 word731 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19670 a_2162_n113516# a_2112_n66# a_1898_n113516# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19671 a_50_n99600# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19672 word71 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19673 word144 A0 a_2294_n20648# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19674 a_1238_n58846# A5 a_974_n58846# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19675 a_2162_n19938# a_2112_n66# a_2030_n19938# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19676 a_2162_n28316# a_2112_n66# a_1898_n28316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19677 word505 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19678 a_1634_n45072# a_1584_n66# a_1370_n45072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19679 word202 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19680 word401 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19681 word474 A0 a_2162_n67508# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19682 a_974_n114794# A6 a_710_n114794# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19683 word410 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19684 a_2162_n97612# a_2112_n66# a_1898_n97612# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19685 word445 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19686 a_1898_n135242# a_1848_n66# a_1766_n135242# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19687 a_1898_n126864# a_1848_n66# a_1634_n126864# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19688 GND A3 word195 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19689 GND A7 word877 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19690 GND A9 word129 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19691 a_2030_n135526# A2 a_1634_n135526# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19692 word36 A0 a_2294_n5312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19693 a_2294_n17950# A1 a_1898_n17950# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19694 a_2294_n26328# A1 a_2030_n26328# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19695 a_314_n129278# a_264_n66# a_50_n129278# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19696 GND A9 word287 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19697 a_2162_n10850# a_2112_n66# a_2030_n10850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19698 word407 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19699 word466 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19700 a_710_n14968# A7 a_446_n14968# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19701 a_1502_n9288# A4 a_1238_n9288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19702 word788 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19703 GND A5 word192 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19704 a_2294_n95624# A1 a_2030_n95624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19705 GND A1 word941 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19706 word468 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19707 a_1634_n74466# a_1584_n66# a_1502_n74466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19708 a_2162_n128426# a_2112_n66# a_1898_n128426# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19709 word717 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19710 a_1634_n124166# a_1584_n66# a_1502_n124166# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19711 a_314_n120190# a_264_n66# a_50_n120190# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19712 a_1106_n123598# a_1056_n66# a_842_n123598# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19713 a_1634_n115788# a_1584_n66# a_1502_n115788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19714 word610 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19715 a_1898_n103292# a_1848_n66# a_1766_n103292# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19716 GND A9 word67 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19717 word178 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19718 a_1502_n87388# A4 a_1106_n87388# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19719 GND A6 word799 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19720 a_578_n105422# a_528_n66# a_446_n105422# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19721 a_2030_n103576# A2 a_1634_n103576# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19722 a_710_n52740# A7 a_314_n52740# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19723 GND A5 word399 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19724 GND A5 word458 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19725 word860 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19726 word995 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19727 word362 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19728 a_1238_n73046# A5 a_974_n73046# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19729 a_1238_n64668# A5 a_842_n64668# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19730 word713 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19731 GND A9 word451 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19732 a_2162_n34138# a_2112_n66# a_1898_n34138# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19733 GND A9 word392 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19734 a_710_n38256# A7 a_314_n38256# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19735 GND A1 word716 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19736 word383 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19737 word984 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19738 word201 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19739 word131 a_2376_n66# a_2162_n18802# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19740 word857 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19741 word781 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19742 a_1898_n132686# a_1848_n66# a_1766_n132686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19743 a_446_n15536# A8 a_182_n15536# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19744 GND A6 word62 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19745 word444 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19746 GND A3 word295 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19747 word763 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19748 GND A9 word170 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19749 a_2030_n141348# A2 a_1766_n141348# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19750 a_2294_n32150# A1 a_2030_n32150# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19751 a_314_n135100# a_264_n66# a_50_n135100# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19752 word669 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19753 a_578_n134816# a_528_n66# a_314_n134816# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19754 word18 A0 a_2162_n2756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19755 a_446_n84832# A8 a_50_n84832# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19756 word507 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19757 GND A5 word665 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19758 word921 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19759 GND A6 word904 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19760 GND A7 word816 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19761 word920 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19762 a_1766_n139360# A3 a_1370_n139360# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19763 GND A1 word824 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19764 GND A1 word765 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19765 a_446_n103008# A8 a_50_n103008# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19766 a_1106_n5454# a_1056_n66# a_974_n5454# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19767 a_710_n76028# A7 a_446_n76028# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19768 a_2030_n58136# A2 a_1634_n58136# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19769 word509 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19770 GND A9 word226 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19771 a_2030_n118486# A2 a_1766_n118486# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19772 word649 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19773 word965 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19774 word927 a_2376_n66# a_2162_n131834# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19775 word290 A0 a_2162_n41380# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19776 word759 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19777 a_2162_n71484# a_2112_n66# a_1898_n71484# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19778 a_446_n102582# A8 a_50_n102582# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19779 a_2294_n78584# A1 a_2030_n78584# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19780 GND A1 word821 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19781 word620 A0 a_2294_n88240# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19782 GND A3 word705 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19783 word1021 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19784 word827 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19785 a_578_n102866# a_528_n66# a_446_n102866# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19786 word549 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19787 word705 a_2376_n66# a_2294_n100310# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19788 word490 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19789 GND A9 word275 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19790 GND A5 word791 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19791 word676 A0 a_2294_n96192# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19792 GND A9 word492 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19793 a_1502_n123314# A4 a_1106_n123314# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19794 a_710_n111528# A7 a_314_n111528# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19795 GND A9 word433 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19796 a_1502_n114936# A4 a_1106_n114936# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19797 a_1106_n15962# a_1056_n66# a_842_n15962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19798 a_710_n44078# A7 a_314_n44078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19799 GND A8 word13 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19800 a_446_n99742# A8 a_50_n99742# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19801 a_1370_n25618# a_1320_n66# a_1106_n25618# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19802 GND A5 word338 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19803 GND A8 word115 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19804 a_2162_n102298# a_2112_n66# a_1898_n102298# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19805 word740 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19806 word231 a_2376_n66# a_2162_n33002# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19807 a_1766_n64810# A3 a_1502_n64810# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19808 word614 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19809 a_2162_n17098# a_2112_n66# a_1898_n17098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19810 word956 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19811 a_446_n21358# A8 a_182_n21358# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19812 GND A1 word108 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19813 GND A6 word44 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19814 a_1370_n94914# a_1320_n66# a_1238_n94914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19815 a_1634_n95198# a_1584_n66# a_1370_n95198# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19816 word695 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19817 a_446_n12980# A8 a_182_n12980# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19818 GND A8 word662 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19819 GND A8 word603 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19820 GND A8 word732 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19821 GND A8 word171 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19822 a_2162_n86394# a_2112_n66# a_1898_n86394# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19823 word745 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19824 a_578_n140638# a_528_n66# a_314_n140638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19825 word63 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19826 a_446_n90654# A8 a_50_n90654# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19827 GND A1 word596 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19828 a_2294_n106558# A1 a_1898_n106558# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19829 GND A6 word945 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19830 GND A1 word865 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19831 a_1238_n112238# A5 a_974_n112238# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19832 a_446_n342# A8 a_182_n342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19833 GND A2 word232 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19834 a_1106_n53734# a_1056_n66# a_842_n53734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19835 a_1106_n62112# a_1056_n66# a_974_n62112# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19836 a_1238_n103860# A5 a_842_n103860# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19837 GND A9 word3 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19838 word508 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19839 a_1238_n85400# A5 a_842_n85400# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19840 GND A5 word896 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19841 a_1502_n138224# A4 a_1238_n138224# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19842 a_1766_n41238# A3 a_1502_n41238# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19843 GND A3 word866 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19844 a_710_n126438# A7 a_314_n126438# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19845 a_2162_n1052# a_2112_n66# a_1898_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19846 a_1766_n32860# A3 a_1502_n32860# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19847 GND A8 word59 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19848 GND A3 word807 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19849 a_1370_n71342# a_1320_n66# a_1106_n71342# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19850 GND A0 word974 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19851 word807 a_2376_n66# a_2162_n114794# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19852 word347 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19853 a_1370_n62964# a_1320_n66# a_1106_n62964# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19854 word277 a_2376_n66# a_2294_n39534# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19855 a_1766_n79720# A3 a_1370_n79720# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19856 a_446_n27890# A8 a_182_n27890# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19857 a_446_n36268# A8 a_182_n36268# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19858 a_1766_n18376# A3 a_1502_n18376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19859 word286 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19860 a_974_n3182# A6 a_710_n3182# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19861 GND A1 word40 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19862 GND A4 word929 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19863 word909 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19864 GND A4 word870 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19865 GND A7 word561 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19866 GND A1 word701 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19867 GND A5 word27 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19868 a_1370_n31440# a_1320_n66# a_1238_n31440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19869 a_2162_n8010# a_2112_n66# a_1898_n8010# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19870 word283 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19871 a_974_n61402# A6 a_578_n61402# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19872 word839 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19873 word213 a_2376_n66# a_2294_n30446# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19874 GND A2 word337 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19875 a_1106_n68644# a_1056_n66# a_842_n68644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19876 a_1238_n118770# A5 a_842_n118770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19877 GND A4 word768 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19878 a_1502_n106274# A4 a_1106_n106274# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19879 word997 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19880 GND A1 word149 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19881 word820 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19882 word543 a_2376_n66# a_2162_n77306# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19883 word554 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19884 word964 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19885 GND A8 word644 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19886 GND A7 word339 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19887 word845 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19888 a_50_n117918# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19889 a_446_n74040# A8 a_50_n74040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19890 GND A1 word420 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19891 GND A0 word462 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19892 GND A7 word280 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19893 GND A8 word714 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19894 a_4084_164# A4 GND GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X19895 GND A1 word637 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19896 word971 a_2376_n66# a_2162_n138082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19897 a_182_n12412# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19898 word45 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19899 a_1370_n86252# a_1320_n66# a_1238_n86252# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19900 GND A7 word14 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19901 a_842_n69922# a_792_n66# a_578_n69922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19902 word775 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19903 GND A8 word542 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19904 GND A6 word179 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19905 word181 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19906 GND A4 word704 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19907 word973 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19908 a_1370_n135384# a_1320_n66# a_1106_n135384# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19909 a_1898_n33712# a_1848_n66# a_1634_n33712# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19910 a_446_n2472# A8 a_182_n2472# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19911 GND A1 word476 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19912 GND A2 word544 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19913 GND A6 word667 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19914 GND A4 word975 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19915 a_1106_n45072# a_1056_n66# a_974_n45072# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19916 a_578_n28742# a_528_n66# a_446_n28742# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19917 GND A4 word174 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19918 GND A7 word605 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19919 a_974_n76312# A6 a_710_n76312# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19920 GND A7 word114 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19921 word259 a_2376_n66# a_2162_n36978# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19922 GND A0 word296 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19923 a_710_n109398# A7 a_314_n109398# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19924 a_182_n41806# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19925 a_314_n48906# a_264_n66# a_182_n48906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19926 a_1502_n23914# A4 a_1106_n23914# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19927 a_446_n9430# A8 a_182_n9430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19928 GND A7 word602 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19929 a_1766_n93494# A3 a_1370_n93494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19930 a_182_n27322# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19931 a_182_n18944# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19932 GND A5 word9 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19933 word880 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19934 a_578_n66514# a_528_n66# a_314_n66514# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19935 GND A4 word809 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19936 a_1898_n48622# a_1848_n66# a_1766_n48622# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19937 GND A6 word442 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19938 GND A4 word750 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19939 a_1238_n768# A5 a_974_n768# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19940 a_50_n88808# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19941 word51 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19942 word654 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19943 GND A5 word4 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19944 GND A5 word983 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19945 GND A0 word790 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19946 a_50_n132118# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19947 GND A7 word380 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19948 word525 a_2376_n66# a_2294_n74750# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19949 GND A0 word562 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19950 a_50_n123740# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19951 a_974_n44362# A6 a_710_n44362# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19952 GND A1 word520 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19953 word31 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19954 word742 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19955 a_842_n84122# a_792_n66# a_710_n84122# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19956 word274 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19957 word222 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19958 word782 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19959 a_50_n109256# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19960 GND A0 word342 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19961 word723 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19962 a_182_n56716# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19963 a_50_n131692# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19964 a_1502_n47202# A4 a_1238_n47202# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19965 word432 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19966 word267 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19967 GND A3 a_1584_n66# GND sky130_fd_pr__nfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X19968 a_578_n95908# a_528_n66# a_446_n95908# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19969 a_314_n140922# a_264_n66# a_50_n140922# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19970 GND A2 word585 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19971 word712 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19972 a_1502_n141490# A4 a_1106_n141490# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19973 GND A5 word919 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19974 GND A2 word784 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19975 a_578_n34564# a_528_n66# a_446_n34564# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19976 a_1898_n16672# a_1848_n66# a_1766_n16672# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19977 a_974_n73756# A6 a_710_n73756# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19978 a_1106_n89376# a_1056_n66# a_842_n89376# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19979 a_182_n7016# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19980 GND A0 word120 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19981 word210 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19982 word359 a_2376_n66# a_2162_n51178# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19983 GND A6 word547 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19984 a_314_n63106# a_264_n66# a_182_n63106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19985 a_50_n100168# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19986 word949 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19987 word1008 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19988 a_314_n54728# a_264_n66# a_182_n54728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19989 word700 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19990 word689 a_2376_n66# a_2294_n98038# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19991 a_50_n138650# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19992 a_974_n59272# A6 a_578_n59272# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19993 GND A0 word608 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19994 a_2030_n5028# A2 a_1766_n5028# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19995 a_842_n52172# a_792_n66# a_710_n52172# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X19996 word639 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19997 GND A0 word176 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X19998 word474 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X19999 word934 A0 a_2162_n132828# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20000 a_182_n33144# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20001 a_1502_n15252# A4 a_1106_n15252# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20002 a_182_n24766# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20003 word386 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20004 a_578_n72336# a_528_n66# a_314_n72336# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20005 a_1106_n80288# a_1056_n66# a_974_n80288# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20006 word887 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20007 a_710_n5170# A7 a_446_n5170# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20008 a_578_n63958# a_528_n66# a_314_n63958# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20009 a_1898_n54444# a_1848_n66# a_1634_n54444# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20010 word537 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20011 word832 A0 a_2294_n118344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20012 a_50_n94630# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20013 word33 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20014 GND A3 word23 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20015 GND A2 word690 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20016 a_842_n12270# a_792_n66# a_710_n12270# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20017 a_974_n19370# A6 a_578_n19370# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20018 word817 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20019 GND A2 word889 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20020 a_1634_n31724# a_1584_n66# a_1370_n31724# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20021 a_1634_n40102# a_1584_n66# a_1370_n40102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20022 word539 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20023 word598 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20024 word758 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20025 GND A4 word320 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20026 word532 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20027 word591 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20028 a_974_n97044# A6 a_578_n97044# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20029 a_50_n106700# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20030 a_50_n115078# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20031 a_182_n62538# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20032 a_314_n69638# a_264_n66# a_182_n69638# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20033 GND A3 word160 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20034 a_314_n124308# a_264_n66# a_50_n124308# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20035 a_1634_n119906# a_1584_n66# a_1502_n119906# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20036 word431 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20037 a_314_n115930# a_264_n66# a_50_n115930# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20038 a_842_n67082# a_792_n66# a_578_n67082# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20039 a_1898_n83838# a_1848_n66# a_1634_n83838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20040 word161 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20041 word1006 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20042 a_1898_n22494# a_1848_n66# a_1634_n22494# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20043 a_1238_n30304# A5 a_842_n30304# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20044 a_842_n120474# a_792_n66# a_710_n120474# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20045 a_182_n39676# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20046 a_182_n48054# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20047 a_1238_n21926# A5 a_974_n21926# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20048 word310 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20049 a_1898_n69354# a_1848_n66# a_1766_n69354# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20050 a_314_n123882# a_264_n66# a_50_n123882# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20051 GND A6 word647 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20052 a_182_n4460# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20053 word141 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20054 a_314_n60550# a_264_n66# a_182_n60550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20055 GND A3 word546 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20056 GND A3 word69 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20057 word331 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20058 a_974_n133112# A6 a_578_n133112# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20059 a_1634_n110818# a_1584_n66# a_1502_n110818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20060 word366 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20061 word725 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20062 a_1502_n82418# A4 a_1238_n82418# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20063 GND A0 word590 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20064 word112 A0 a_2294_n16104# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20065 word888 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20066 VDD A0 a_2376_n66# VDD sky130_fd_pr__pfet_01v8 ad=0.1548 pd=1.58 as=0.1548 ps=1.58 w=0.43 l=0.17
X20067 a_314_n37688# a_264_n66# a_182_n37688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20068 a_314_n46066# a_264_n66# a_182_n46066# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20069 GND A4 word583 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20070 GND A4 word642 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20071 a_182_n30588# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20072 GND A3 word324 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20073 a_1898_n51888# a_1848_n66# a_1634_n51888# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20074 a_1898_n60266# a_1848_n66# a_1766_n60266# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20075 GND A0 word488 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20076 a_1502_n59556# A4 a_1106_n59556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20077 a_314_n139218# a_264_n66# a_50_n139218# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20078 word698 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20079 word814 A0 a_2162_n115788# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20080 a_1502_n81992# A4 a_1238_n81992# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20081 word47 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20082 word85 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20083 a_1634_n15110# a_1584_n66# a_1502_n15110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20084 a_1898_n98748# a_1848_n66# a_1766_n98748# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20085 word858 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20086 GND A2 word930 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20087 GND A5 word262 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20088 word207 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20089 word580 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20090 word799 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20091 a_1238_n36836# A5 a_974_n36836# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20092 a_578_n55296# a_528_n66# a_314_n55296# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20093 a_50_n77590# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20094 word415 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20095 GND A3 word321 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20096 a_974_n94488# A6 a_578_n94488# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20097 word573 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20098 word106 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20099 a_314_n138792# a_264_n66# a_50_n138792# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20100 GND A2 word769 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20101 word187 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20102 word255 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20103 a_1502_n50468# A4 a_1106_n50468# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20104 a_314_n130130# a_264_n66# a_50_n130130# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20105 a_1634_n134106# a_1584_n66# a_1502_n134106# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20106 a_1106_n133538# a_1056_n66# a_974_n133538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20107 GND A4 word200 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20108 a_2162_n75602# a_2112_n66# a_2030_n75602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20109 word290 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20110 a_1898_n113232# a_1848_n66# a_1634_n113232# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20111 word471 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20112 word830 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20113 word248 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20114 a_1502_n97328# A4 a_1106_n97328# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20115 word988 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20116 GND A7 word781 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20117 a_182_n45498# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20118 GND A3 word99 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20119 word473 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20120 word311 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20121 a_578_n93068# a_528_n66# a_446_n93068# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20122 word414 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20123 a_1898_n66798# a_1848_n66# a_1766_n66798# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20124 a_1238_n74608# A5 a_974_n74608# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20125 word978 A0 a_2162_n139076# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20126 GND A9 word462 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20127 a_1238_n13264# A5 a_842_n13264# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20128 word190 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20129 word372 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20130 a_2294_n73614# A1 a_1898_n73614# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20131 a_1766_n200# A3 a_1502_n200# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20132 a_710_n39818# A7 a_314_n39818# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20133 word904 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20134 a_974_n130556# A6 a_578_n130556# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20135 GND A7 word0 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20136 word453 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20137 word685 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20138 word986 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20139 word94 A0 a_2162_n13548# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20140 a_1634_n102156# a_1584_n66# a_1502_n102156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20141 word678 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20142 a_1634_n99316# a_1584_n66# a_1370_n99316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20143 a_974_n116072# A6 a_710_n116072# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20144 a_2162_n43652# a_2112_n66# a_2030_n43652# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20145 a_1634_n29594# a_1584_n66# a_1502_n29594# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20146 GND A6 word703 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20147 a_1502_n65378# A4 a_1238_n65378# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20148 a_314_n145040# a_264_n66# a_50_n145040# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20149 word582 A0 a_2162_n82844# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20150 a_1766_n102440# A3 a_1370_n102440# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20151 word680 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20152 word395 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20153 word991 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20154 a_1898_n128142# a_1848_n66# a_1766_n128142# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20155 word766 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20156 word518 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20157 a_2030_n12838# A2 a_1634_n12838# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20158 word705 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20159 word511 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20160 GND A7 word827 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20161 GND A7 word886 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20162 word579 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20163 GND A9 word296 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20164 a_1634_n90228# a_1584_n66# a_1370_n90228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20165 GND A9 word237 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20166 a_710_n16246# A7 a_446_n16246# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20167 word88 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20168 a_2294_n41664# A1 a_1898_n41664# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20169 a_578_n99600# a_528_n66# a_446_n99600# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20170 a_1634_n81850# a_1584_n66# a_1370_n81850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20171 a_2162_n135810# a_2112_n66# a_2030_n135810# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20172 word360 A0 a_2294_n51320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20173 a_1238_n28174# A5 a_842_n28174# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20174 GND A3 word692 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20175 a_1634_n131550# a_1584_n66# a_1370_n131550# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20176 a_1238_n19796# A5 a_974_n19796# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20177 GND A3 word836 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20178 word230 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20179 word289 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20180 a_1634_n58988# a_1584_n66# a_1370_n58988# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20181 a_1634_n67366# a_1584_n66# a_1370_n67366# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20182 a_710_n85542# A7 a_446_n85542# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20183 word576 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20184 a_2162_n143762# a_2112_n66# a_2030_n143762# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20185 a_314_n113090# a_264_n66# a_50_n113090# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20186 a_1106_n116498# a_1056_n66# a_974_n116498# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20187 word135 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20188 a_2030_n50610# A2 a_1766_n50610# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20189 a_2162_n58562# a_2112_n66# a_2030_n58562# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20190 word560 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20191 a_1634_n108688# a_1584_n66# a_1370_n108688# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20192 GND A5 word78 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20193 GND A9 word503 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20194 a_1106_n25902# a_1056_n66# a_974_n25902# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20195 a_710_n54018# A7 a_314_n54018# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20196 word623 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20197 word682 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20198 a_2030_n27748# A2 a_1766_n27748# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20199 a_710_n45640# A7 a_314_n45640# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20200 GND A5 word408 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20201 GND A8 word24 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20202 word354 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20203 word945 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20204 GND A9 word71 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20205 word312 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20206 GND A5 word349 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20207 word435 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20208 a_1238_n57568# A5 a_974_n57568# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20209 word616 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20210 a_2162_n103860# a_2112_n66# a_2030_n103860# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20211 word625 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20212 GND A9 word401 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20213 GND A9 word342 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20214 a_2162_n18660# a_2112_n66# a_2030_n18660# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20215 a_2294_n56574# A1 a_1898_n56574# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20216 a_1634_n96760# a_1584_n66# a_1502_n96760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20217 a_446_n22920# A8 a_182_n22920# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20218 a_710_n53592# A7 a_314_n53592# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20219 word333 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20220 GND A8 word241 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20221 GND A8 word743 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20222 word866 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20223 word815 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20224 a_2162_n87956# a_2112_n66# a_2030_n87956# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20225 word731 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20226 a_1766_n82702# A3 a_1502_n82702# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20227 GND A7 word43 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20228 GND A5 word285 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20229 a_446_n30872# A8 a_182_n30872# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20230 GND A7 word868 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20231 GND A9 word120 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20232 GND A2 word243 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20233 a_1502_n101304# A4 a_1238_n101304# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20234 a_1370_n139502# a_1320_n66# a_1238_n139502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20235 a_2030_n134248# A2 a_1766_n134248# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20236 a_578_n127716# a_528_n66# a_314_n127716# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20237 word871 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20238 a_446_n77732# A8 a_50_n77732# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20239 a_1238_n95340# A5 a_974_n95340# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20240 a_710_n13690# A7 a_446_n13690# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20241 word929 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20242 a_2294_n85968# A1 a_1898_n85968# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20243 word459 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20244 GND A9 word176 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20245 GND A1 word932 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20246 a_1238_n121752# A5 a_842_n121752# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20247 word599 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20248 word801 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20249 word877 a_2376_n66# a_2294_n124734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20250 a_710_n82986# A7 a_446_n82986# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20251 GND A5 word671 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20252 a_2162_n127148# a_2112_n66# a_1898_n127148# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20253 a_2162_n118770# a_2112_n66# a_2030_n118770# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20254 word240 A0 a_2294_n34280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20255 word926 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20256 a_1370_n130414# a_1320_n66# a_1238_n130414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20257 a_1766_n28316# A3 a_1502_n28316# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20258 GND A7 word301 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20259 a_974_n4744# A6 a_710_n4744# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20260 a_1766_n50752# A3 a_1502_n50752# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20261 GND A1 word441 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20262 GND A9 word58 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20263 word169 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20264 word979 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20265 GND A6 word790 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20266 GND A7 word631 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20267 word971 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20268 a_578_n104144# a_528_n66# a_446_n104144# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20269 a_1370_n107552# a_1320_n66# a_1106_n107552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20270 a_2030_n33570# A2 a_1634_n33570# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20271 GND A5 word390 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20272 word626 A0 a_2162_n89092# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20273 word704 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20274 a_1238_n128710# A5 a_974_n128710# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20275 GND A7 word79 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20276 GND A9 word383 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20277 GND A3 word711 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20278 GND A4 word996 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20279 GND A1 word160 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20280 word711 a_2376_n66# a_2162_n101162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20281 word975 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20282 word915 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20283 a_1370_n40954# a_1320_n66# a_1238_n40954# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20284 a_1766_n57710# A3 a_1370_n57710# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20285 GND A8 word223 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20286 a_2162_n93778# a_2112_n66# a_2030_n93778# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20287 word713 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20288 GND A7 word567 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20289 word906 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20290 GND A3 word982 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20291 a_1238_n136662# A5 a_842_n136662# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20292 a_2294_n122320# A1 a_1898_n122320# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20293 a_1634_n88098# a_1584_n66# a_1502_n88098# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20294 a_446_n14258# A8 a_182_n14258# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20295 GND A7 word76 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20296 GND A8 word612 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20297 GND A1 word216 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20298 GND A7 word25 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20299 GND A8 word553 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20300 word946 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20301 GND A4 word715 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20302 GND A7 word850 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20303 word984 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20304 a_1370_n145324# a_1320_n66# a_1106_n145324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20305 a_2030_n140070# A2 a_1634_n140070# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20306 GND A4 word774 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20307 a_578_n133538# a_528_n66# a_314_n133538# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20308 GND A8 word121 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20309 a_446_n83554# A8 a_50_n83554# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20310 a_2294_n130272# A1 a_1898_n130272# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20311 a_2294_n121894# A1 a_2030_n121894# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20312 GND A2 word123 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20313 word500 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20314 a_2294_n91790# A1 a_1898_n91790# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20315 GND A3 word918 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20316 word458 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20317 word724 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20318 word399 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20319 a_1634_n4602# a_1584_n66# a_1370_n4602# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20320 GND A7 word125 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20321 word329 a_2376_n66# a_2294_n46918# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20322 word750 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20323 GND A9 word488 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20324 word920 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20325 a_710_n119338# A7 a_314_n119338# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20326 GND A1 word265 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20327 GND A1 word324 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20328 GND A2 word611 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20329 GND A3 word816 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20330 GND A3 word757 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20331 a_1766_n25760# A3 a_1370_n25760# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20332 word757 a_2376_n66# a_2294_n107694# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20333 GND A9 word40 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20334 a_1106_n15110# a_1056_n66# a_842_n15110# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20335 a_842_n47912# a_792_n66# a_710_n47912# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20336 word721 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20337 a_2294_n137230# A1 a_1898_n137230# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20338 a_1370_n113374# a_1320_n66# a_1238_n113374# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20339 a_446_n29168# A8 a_182_n29168# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20340 a_578_n101588# a_528_n66# a_446_n101588# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20341 GND A1 word49 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20342 GND A1 word321 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20343 GND A4 word879 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20344 GND A5 word782 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20345 GND A6 word512 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20346 a_710_n110250# A7 a_314_n110250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20347 GND A5 word723 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20348 a_1106_n14684# a_1056_n66# a_842_n14684# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20349 a_1106_n23062# a_1056_n66# a_974_n23062# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20350 a_446_n98464# A8 a_50_n98464# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20351 word665 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20352 a_2294_n145182# A1 a_1898_n145182# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20353 GND A0 word860 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20354 word233 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20355 word163 a_2376_n66# a_2162_n23346# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20356 word947 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20357 word1006 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20358 a_446_n20080# A8 a_182_n20080# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20359 GND A0 word82 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20360 word1023 a_2376_n66# a_2162_n145466# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20361 GND A4 word876 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20362 word812 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20363 GND A6 word35 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20364 a_1370_n93636# a_1320_n66# a_1238_n93636# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20365 a_710_n8862# A7 a_446_n8862# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20366 word987 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20367 GND A8 word594 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20368 GND A0 word412 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20369 word651 a_2376_n66# a_2162_n92642# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20370 GND A0 word916 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20371 word795 a_3028_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20372 a_842_n15962# a_792_n66# a_710_n15962# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20373 a_50_n141632# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20374 a_2294_n105280# A1 a_1898_n105280# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20375 word25 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20376 a_446_n80998# A8 a_50_n80998# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20377 a_1766_n71484# A3 a_1370_n71484# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20378 GND A5 word989 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20379 GND A6 word129 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20380 word131 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20381 word826 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20382 a_1106_n52456# a_1056_n66# a_842_n52456# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20383 GND A6 word287 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20384 word341 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20385 word429 a_2376_n66# a_2294_n61118# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20386 word440 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20387 a_1106_n99316# a_1056_n66# a_974_n99316# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20388 a_50_n110108# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20389 a_1502_n128568# A4 a_1238_n128568# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20390 a_710_n125160# A7 a_314_n125160# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20391 a_50_n101730# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20392 a_974_n22352# A6 a_578_n22352# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20393 GND A1 word365 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20394 a_1370_n39250# a_1320_n66# a_1238_n39250# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20395 GND A8 word50 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20396 GND A7 word555 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20397 a_842_n53734# a_792_n66# a_710_n53734# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20398 a_1370_n61686# a_1320_n66# a_1106_n61686# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20399 word209 a_2376_n66# a_2294_n29878# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20400 GND A0 word246 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20401 word859 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20402 a_1766_n17098# A3 a_1370_n17098# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20403 GND A1 word204 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20404 a_182_n34706# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20405 GND A8 word699 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20406 a_1106_n81850# a_1056_n66# a_974_n81850# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20407 a_1106_n90228# a_1056_n66# a_842_n90228# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20408 word898 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20409 GND A1 word692 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20410 word751 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20411 GND A7 word552 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20412 word116 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20413 a_974_n60124# A6 a_578_n60124# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20414 word830 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20415 word145 a_2376_n66# a_2294_n20790# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20416 a_578_n59414# a_528_n66# a_314_n59414# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20417 GND A6 word392 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20418 word988 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20419 a_842_n139502# a_792_n66# a_578_n139502# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20420 GND A1 word140 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20421 a_974_n98606# A6 a_578_n98606# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20422 word475 a_2376_n66# a_2162_n67650# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20423 GND A7 word330 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20424 GND A0 word740 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20425 GND A8 word635 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20426 a_50_n116640# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20427 a_50_n125018# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20428 a_842_n30162# a_792_n66# a_578_n30162# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20429 a_974_n37262# A6 a_710_n37262# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20430 a_1766_n1052# A3 a_1502_n1052# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20431 word111 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20432 GND A1 word569 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20433 a_182_n11134# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20434 word12 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20435 a_1370_n76596# a_1320_n66# a_1238_n76596# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20436 GND A6 word170 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20437 a_842_n68644# a_792_n66# a_578_n68644# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20438 word172 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20439 word231 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20440 word382 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20441 a_446_n1194# A8 a_182_n1194# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20442 a_182_n49616# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20443 a_50_n124592# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20444 a_1898_n6874# a_1848_n66# a_1634_n6874# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20445 a_314_n133822# a_264_n66# a_50_n133822# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20446 a_1106_n96760# a_1056_n66# a_974_n96760# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20447 GND A6 word658 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20448 GND A4 word224 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20449 a_578_n27464# a_528_n66# a_446_n27464# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20450 word27 a_3820_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20451 GND A4 word165 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20452 a_842_n107552# a_792_n66# a_578_n107552# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20453 word65 a_2376_n66# a_2294_n9430# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20454 GND A5 word64 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20455 a_974_n75034# A6 a_710_n75034# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20456 a_50_n80572# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20457 a_1766_n8010# A3 a_1370_n8010# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20458 word309 a_2376_n66# a_2294_n44078# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20459 word436 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20460 GND A6 word556 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20461 GND A0 word660 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20462 a_2294_n3182# A1 a_1898_n3182# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20463 word958 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20464 a_314_n56006# a_264_n66# a_182_n56006# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20465 GND A0 word228 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20466 GND A4 word653 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20467 a_182_n40528# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20468 a_314_n47628# a_264_n66# a_182_n47628# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20469 GND A2 word17 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20470 a_1106_n105706# a_1056_n66# a_842_n105706# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20471 GND A4 word68 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20472 a_1898_n70206# a_1848_n66# a_1634_n70206# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20473 GND A0 word558 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20474 word939 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20475 word884 A0 a_2294_n125728# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20476 a_1766_n7584# A3 a_1370_n7584# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20477 GND A0 word126 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20478 GND A4 word551 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20479 a_1502_n91932# A4 a_1238_n91932# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20480 a_182_n17666# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20481 a_182_n26044# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20482 word157 a_4084_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20483 GND A6 word275 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20484 a_578_n65236# a_528_n66# a_314_n65236# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20485 a_1898_n47344# a_1848_n66# a_1634_n47344# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20486 GND A6 word433 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20487 a_842_n145324# a_792_n66# a_578_n145324# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20488 a_842_n136946# a_792_n66# a_578_n136946# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20489 a_50_n87530# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20490 word42 a_4348_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20491 a_578_n56858# a_528_n66# a_314_n56858# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20492 GND A3 word391 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20493 a_974_n111102# A6 a_710_n111102# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20494 word117 a_4612_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20495 a_974_n43084# A6 a_710_n43084# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20496 GND A0 word494 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20497 word548 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20498 word767 a_5404_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20499 word421 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20500 a_1634_n24624# a_1584_n66# a_1502_n24624# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20501 a_1502_n60408# A4 a_1106_n60408# VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20502 word22 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20503 GND A4 word270 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20504 word360 a_5140_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20505 GND A4 word428 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20506 word541 a_3556_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20507 a_50_n95482# a_0_n66# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20508 GND A4 word1 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20509 word213 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20510 a_1634_n8294# a_1584_n66# a_1370_n8294# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20511 word714 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20512 a_182_n55438# A9 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20513 word718 A0 a_2162_n102156# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20514 a_1502_n37546# A4 a_1238_n37546# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20515 a_314_n117208# a_264_n66# a_50_n117208# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20516 word322 a_3292_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.10535 pd=0.92 as=0.1763 ps=1.68 w=0.43 l=0.17
X20517 GND A4 word326 GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
X20518 a_1898_n85116# a_1848_n66# a_1766_n85116# VDD sky130_fd_pr__pfet_01v8 ad=0.1763 pd=1.68 as=0.10535 ps=0.92 w=0.43 l=0.17
X20519 word484 a_4876_164# GND GND sky130_fd_pr__nfet_01v8 ad=0.1763 pd=1.68 as=0.1763 ps=1.68 w=0.43 l=0.17
.ends

.subckt counter_4 CLK Q0 Q1 Q2 Q3 GND VDD
Xtff_0 tff_0/T CLK inv_1/Y Q2 tff_0/~Q GND VDD tff
Xtff_1 VDD CLK inv_1/Y Q0 tff_1/~Q GND VDD tff
Xtff_2 tff_2/T CLK inv_1/Y Q1 tff_2/~Q GND VDD tff
Xtff_3 tff_3/T CLK inv_1/Y Q3 tff_3/~Q GND VDD tff
Xinv_1 VDD GND CLK inv_1/Y inv
Xinv_2 VDD GND inv_2/A tff_2/T inv
Xinv_3 VDD GND inv_3/A tff_0/T inv
Xinv_4 VDD GND inv_4/A tff_3/T inv
Xnand_0 VDD GND tff_0/T inv_4/A Q2 nand
Xnand_1 VDD GND VDD inv_2/A Q0 nand
Xnand_2 VDD GND tff_2/T inv_3/A Q1 nand
.ends

*.subckt func_gen_8_connected CLK Freq0 Freq1 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 Wave0 Wave1
Xmemory_8_0 memory_8_0/word0 memory_8_0/word1 memory_8_0/word2 memory_8_0/word3 memory_8_0/word4
+ memory_8_0/word5 memory_8_0/word6 memory_8_0/word7 memory_8_0/word8 memory_8_0/word9
+ memory_8_0/word10 memory_8_0/word11 memory_8_0/word12 memory_8_0/word13 memory_8_0/word14
+ memory_8_0/word15 memory_8_0/word16 memory_8_0/word17 memory_8_0/word18 memory_8_0/word19
+ memory_8_0/word20 memory_8_0/word21 memory_8_0/word22 memory_8_0/word23 memory_8_0/word24
+ memory_8_0/word25 memory_8_0/word26 memory_8_0/word27 memory_8_0/word28 memory_8_0/word29
+ memory_8_0/word30 memory_8_0/word31 memory_8_0/word32 memory_8_0/word33 memory_8_0/word34
+ memory_8_0/word35 memory_8_0/word36 memory_8_0/word37 memory_8_0/word38 memory_8_0/word39
+ memory_8_0/word40 memory_8_0/word41 memory_8_0/word42 memory_8_0/word43 memory_8_0/word44
+ memory_8_0/word45 memory_8_0/word46 memory_8_0/word47 memory_8_0/word48 memory_8_0/word49
+ memory_8_0/word50 memory_8_0/word51 memory_8_0/word52 memory_8_0/word53 memory_8_0/word54
+ memory_8_0/word55 memory_8_0/word56 memory_8_0/word57 memory_8_0/word58 memory_8_0/word59
+ memory_8_0/word60 memory_8_0/word61 memory_8_0/word62 memory_8_0/word63 memory_8_0/word64
+ memory_8_0/word65 memory_8_0/word66 memory_8_0/word67 memory_8_0/word68 memory_8_0/word69
+ memory_8_0/word70 memory_8_0/word71 memory_8_0/word72 memory_8_0/word73 memory_8_0/word74
+ memory_8_0/word75 memory_8_0/word76 memory_8_0/word77 memory_8_0/word78 memory_8_0/word79
+ memory_8_0/word80 memory_8_0/word81 memory_8_0/word82 memory_8_0/word83 memory_8_0/word84
+ memory_8_0/word85 memory_8_0/word86 memory_8_0/word87 memory_8_0/word88 memory_8_0/word89
+ memory_8_0/word90 memory_8_0/word91 memory_8_0/word92 memory_8_0/word93 memory_8_0/word94
+ memory_8_0/word95 memory_8_0/word96 memory_8_0/word97 memory_8_0/word98 memory_8_0/word99
+ memory_8_0/word100 memory_8_0/word101 memory_8_0/word102 memory_8_0/word103 memory_8_0/word104
+ memory_8_0/word105 memory_8_0/word106 memory_8_0/word107 memory_8_0/word108 memory_8_0/word109
+ memory_8_0/word110 memory_8_0/word111 memory_8_0/word112 memory_8_0/word113 memory_8_0/word114
+ memory_8_0/word115 memory_8_0/word116 memory_8_0/word117 memory_8_0/word118 memory_8_0/word119
+ memory_8_0/word120 memory_8_0/word121 memory_8_0/word122 memory_8_0/word123 memory_8_0/word124
+ memory_8_0/word125 memory_8_0/word126 memory_8_0/word127 memory_8_0/word128 memory_8_0/word129
+ memory_8_0/word130 memory_8_0/word131 memory_8_0/word132 memory_8_0/word133 memory_8_0/word134
+ memory_8_0/word135 memory_8_0/word136 memory_8_0/word137 memory_8_0/word138 memory_8_0/word139
+ memory_8_0/word140 memory_8_0/word141 memory_8_0/word142 memory_8_0/word143 memory_8_0/word144
+ memory_8_0/word145 memory_8_0/word146 memory_8_0/word147 memory_8_0/word148 memory_8_0/word149
+ memory_8_0/word150 memory_8_0/word151 memory_8_0/word152 memory_8_0/word153 memory_8_0/word154
+ memory_8_0/word155 memory_8_0/word156 memory_8_0/word157 memory_8_0/word158 memory_8_0/word159
+ memory_8_0/word160 memory_8_0/word161 memory_8_0/word162 memory_8_0/word163 memory_8_0/word164
+ memory_8_0/word165 memory_8_0/word166 memory_8_0/word167 memory_8_0/word168 memory_8_0/word169
+ memory_8_0/word170 memory_8_0/word171 memory_8_0/word172 memory_8_0/word173 memory_8_0/word174
+ memory_8_0/word175 memory_8_0/word176 memory_8_0/word177 memory_8_0/word178 memory_8_0/word179
+ memory_8_0/word180 memory_8_0/word181 memory_8_0/word182 memory_8_0/word183 memory_8_0/word184
+ memory_8_0/word185 memory_8_0/word186 memory_8_0/word187 memory_8_0/word188 memory_8_0/word189
+ memory_8_0/word190 memory_8_0/word191 memory_8_0/word192 memory_8_0/word193 memory_8_0/word194
+ memory_8_0/word195 memory_8_0/word196 memory_8_0/word197 memory_8_0/word198 memory_8_0/word199
+ memory_8_0/word200 memory_8_0/word201 memory_8_0/word202 memory_8_0/word203 memory_8_0/word204
+ memory_8_0/word205 memory_8_0/word206 memory_8_0/word207 memory_8_0/word208 memory_8_0/word209
+ memory_8_0/word210 memory_8_0/word211 memory_8_0/word212 memory_8_0/word213 memory_8_0/word214
+ memory_8_0/word215 memory_8_0/word216 memory_8_0/word217 memory_8_0/word218 memory_8_0/word219
+ memory_8_0/word220 memory_8_0/word221 memory_8_0/word222 memory_8_0/word223 memory_8_0/word224
+ memory_8_0/word225 memory_8_0/word226 memory_8_0/word227 memory_8_0/word228 memory_8_0/word229
+ memory_8_0/word230 memory_8_0/word231 memory_8_0/word232 memory_8_0/word233 memory_8_0/word234
+ memory_8_0/word235 memory_8_0/word236 memory_8_0/word237 memory_8_0/word238 memory_8_0/word239
+ memory_8_0/word240 memory_8_0/word241 memory_8_0/word242 memory_8_0/word243 memory_8_0/word244
+ memory_8_0/word245 memory_8_0/word246 memory_8_0/word247 memory_8_0/word248 memory_8_0/word249
+ memory_8_0/word250 memory_8_0/word251 memory_8_0/word252 memory_8_0/word253 memory_8_0/word254
+ memory_8_0/word255 memory_8_0/word256 memory_8_0/word257 memory_8_0/word258 memory_8_0/word259
+ memory_8_0/word260 memory_8_0/word261 memory_8_0/word262 memory_8_0/word263 memory_8_0/word264
+ memory_8_0/word265 memory_8_0/word266 memory_8_0/word267 memory_8_0/word268 memory_8_0/word269
+ memory_8_0/word270 memory_8_0/word271 memory_8_0/word272 memory_8_0/word273 memory_8_0/word274
+ memory_8_0/word275 memory_8_0/word276 memory_8_0/word277 memory_8_0/word278 memory_8_0/word279
+ memory_8_0/word280 memory_8_0/word281 memory_8_0/word282 memory_8_0/word283 memory_8_0/word284
+ memory_8_0/word285 memory_8_0/word286 memory_8_0/word287 memory_8_0/word288 memory_8_0/word289
+ memory_8_0/word290 memory_8_0/word291 memory_8_0/word292 memory_8_0/word293 memory_8_0/word294
+ memory_8_0/word295 memory_8_0/word296 memory_8_0/word297 memory_8_0/word298 memory_8_0/word299
+ memory_8_0/word300 memory_8_0/word301 memory_8_0/word302 memory_8_0/word303 memory_8_0/word304
+ memory_8_0/word305 memory_8_0/word306 memory_8_0/word307 memory_8_0/word308 memory_8_0/word309
+ memory_8_0/word310 memory_8_0/word311 memory_8_0/word312 memory_8_0/word313 memory_8_0/word314
+ memory_8_0/word315 memory_8_0/word316 memory_8_0/word317 memory_8_0/word318 memory_8_0/word319
+ memory_8_0/word320 memory_8_0/word321 memory_8_0/word322 memory_8_0/word323 memory_8_0/word324
+ memory_8_0/word325 memory_8_0/word326 memory_8_0/word327 memory_8_0/word328 memory_8_0/word329
+ memory_8_0/word330 memory_8_0/word331 memory_8_0/word332 memory_8_0/word333 memory_8_0/word334
+ memory_8_0/word335 memory_8_0/word336 memory_8_0/word337 memory_8_0/word338 memory_8_0/word339
+ memory_8_0/word340 memory_8_0/word341 memory_8_0/word342 memory_8_0/word343 memory_8_0/word344
+ memory_8_0/word345 memory_8_0/word346 memory_8_0/word347 memory_8_0/word348 memory_8_0/word349
+ memory_8_0/word350 memory_8_0/word351 memory_8_0/word352 memory_8_0/word353 memory_8_0/word354
+ memory_8_0/word355 memory_8_0/word356 memory_8_0/word357 memory_8_0/word358 memory_8_0/word359
+ memory_8_0/word360 memory_8_0/word361 memory_8_0/word362 memory_8_0/word363 memory_8_0/word364
+ memory_8_0/word365 memory_8_0/word366 memory_8_0/word367 memory_8_0/word368 memory_8_0/word369
+ memory_8_0/word370 memory_8_0/word371 memory_8_0/word372 memory_8_0/word373 memory_8_0/word374
+ memory_8_0/word375 memory_8_0/word376 memory_8_0/word377 memory_8_0/word378 memory_8_0/word379
+ memory_8_0/word380 memory_8_0/word381 memory_8_0/word382 memory_8_0/word383 memory_8_0/word384
+ memory_8_0/word385 memory_8_0/word386 memory_8_0/word387 memory_8_0/word388 memory_8_0/word389
+ memory_8_0/word390 memory_8_0/word391 memory_8_0/word392 memory_8_0/word393 memory_8_0/word394
+ memory_8_0/word395 memory_8_0/word396 memory_8_0/word397 memory_8_0/word398 memory_8_0/word399
+ memory_8_0/word400 memory_8_0/word401 memory_8_0/word402 memory_8_0/word403 memory_8_0/word404
+ memory_8_0/word405 memory_8_0/word406 memory_8_0/word407 memory_8_0/word408 memory_8_0/word409
+ memory_8_0/word410 memory_8_0/word411 memory_8_0/word412 memory_8_0/word413 memory_8_0/word414
+ memory_8_0/word415 memory_8_0/word416 memory_8_0/word417 memory_8_0/word418 memory_8_0/word419
+ memory_8_0/word420 memory_8_0/word421 memory_8_0/word422 memory_8_0/word423 memory_8_0/word424
+ memory_8_0/word425 memory_8_0/word426 memory_8_0/word427 memory_8_0/word428 memory_8_0/word429
+ memory_8_0/word430 memory_8_0/word431 memory_8_0/word432 memory_8_0/word433 memory_8_0/word434
+ memory_8_0/word435 memory_8_0/word436 memory_8_0/word437 memory_8_0/word438 memory_8_0/word439
+ memory_8_0/word440 memory_8_0/word441 memory_8_0/word442 memory_8_0/word443 memory_8_0/word444
+ memory_8_0/word445 memory_8_0/word446 memory_8_0/word447 memory_8_0/word448 memory_8_0/word449
+ memory_8_0/word450 memory_8_0/word451 memory_8_0/word452 memory_8_0/word453 memory_8_0/word454
+ memory_8_0/word455 memory_8_0/word456 memory_8_0/word457 memory_8_0/word458 memory_8_0/word459
+ memory_8_0/word460 memory_8_0/word461 memory_8_0/word462 memory_8_0/word463 memory_8_0/word464
+ memory_8_0/word465 memory_8_0/word466 memory_8_0/word467 memory_8_0/word468 memory_8_0/word469
+ memory_8_0/word470 memory_8_0/word471 memory_8_0/word472 memory_8_0/word473 memory_8_0/word474
+ memory_8_0/word475 memory_8_0/word476 memory_8_0/word477 memory_8_0/word478 memory_8_0/word479
+ memory_8_0/word480 memory_8_0/word481 memory_8_0/word482 memory_8_0/word483 memory_8_0/word484
+ memory_8_0/word485 memory_8_0/word486 memory_8_0/word487 memory_8_0/word488 memory_8_0/word489
+ memory_8_0/word490 memory_8_0/word491 memory_8_0/word492 memory_8_0/word493 memory_8_0/word494
+ memory_8_0/word495 memory_8_0/word496 memory_8_0/word497 memory_8_0/word498 memory_8_0/word499
+ memory_8_0/word500 memory_8_0/word501 memory_8_0/word502 memory_8_0/word503 memory_8_0/word504
+ memory_8_0/word505 memory_8_0/word506 memory_8_0/word507 memory_8_0/word508 memory_8_0/word509
+ memory_8_0/word510 memory_8_0/word511 memory_8_0/word512 memory_8_0/word513 memory_8_0/word514
+ memory_8_0/word515 memory_8_0/word516 memory_8_0/word517 memory_8_0/word518 memory_8_0/word519
+ memory_8_0/word520 memory_8_0/word521 memory_8_0/word522 memory_8_0/word523 memory_8_0/word524
+ memory_8_0/word525 memory_8_0/word526 memory_8_0/word527 memory_8_0/word528 memory_8_0/word529
+ memory_8_0/word530 memory_8_0/word531 memory_8_0/word532 memory_8_0/word533 memory_8_0/word534
+ memory_8_0/word535 memory_8_0/word536 memory_8_0/word537 memory_8_0/word538 memory_8_0/word539
+ memory_8_0/word540 memory_8_0/word541 memory_8_0/word542 memory_8_0/word543 memory_8_0/word544
+ memory_8_0/word545 memory_8_0/word546 memory_8_0/word547 memory_8_0/word548 memory_8_0/word549
+ memory_8_0/word550 memory_8_0/word551 memory_8_0/word552 memory_8_0/word553 memory_8_0/word554
+ memory_8_0/word555 memory_8_0/word556 memory_8_0/word557 memory_8_0/word558 memory_8_0/word559
+ memory_8_0/word560 memory_8_0/word561 memory_8_0/word562 memory_8_0/word563 memory_8_0/word564
+ memory_8_0/word565 memory_8_0/word566 memory_8_0/word567 memory_8_0/word568 memory_8_0/word569
+ memory_8_0/word570 memory_8_0/word571 memory_8_0/word572 memory_8_0/word573 memory_8_0/word574
+ memory_8_0/word575 memory_8_0/word576 memory_8_0/word577 memory_8_0/word578 memory_8_0/word579
+ memory_8_0/word580 memory_8_0/word581 memory_8_0/word582 memory_8_0/word583 memory_8_0/word584
+ memory_8_0/word585 memory_8_0/word586 memory_8_0/word587 memory_8_0/word588 memory_8_0/word589
+ memory_8_0/word590 memory_8_0/word591 memory_8_0/word592 memory_8_0/word593 memory_8_0/word594
+ memory_8_0/word595 memory_8_0/word596 memory_8_0/word597 memory_8_0/word598 memory_8_0/word599
+ memory_8_0/word600 memory_8_0/word601 memory_8_0/word602 memory_8_0/word603 memory_8_0/word604
+ memory_8_0/word605 memory_8_0/word606 memory_8_0/word607 memory_8_0/word608 memory_8_0/word609
+ memory_8_0/word610 memory_8_0/word611 memory_8_0/word612 memory_8_0/word613 memory_8_0/word614
+ memory_8_0/word615 memory_8_0/word616 memory_8_0/word617 memory_8_0/word618 memory_8_0/word619
+ memory_8_0/word620 memory_8_0/word621 memory_8_0/word622 memory_8_0/word623 memory_8_0/word624
+ memory_8_0/word625 memory_8_0/word626 memory_8_0/word627 memory_8_0/word628 memory_8_0/word629
+ memory_8_0/word630 memory_8_0/word631 memory_8_0/word632 memory_8_0/word633 memory_8_0/word634
+ memory_8_0/word635 memory_8_0/word636 memory_8_0/word637 memory_8_0/word638 memory_8_0/word639
+ memory_8_0/word640 memory_8_0/word641 memory_8_0/word642 memory_8_0/word643 memory_8_0/word644
+ memory_8_0/word645 memory_8_0/word646 memory_8_0/word647 memory_8_0/word648 memory_8_0/word649
+ memory_8_0/word650 memory_8_0/word651 memory_8_0/word652 memory_8_0/word653 memory_8_0/word654
+ memory_8_0/word655 memory_8_0/word656 memory_8_0/word657 memory_8_0/word658 memory_8_0/word659
+ memory_8_0/word660 memory_8_0/word661 memory_8_0/word662 memory_8_0/word663 memory_8_0/word664
+ memory_8_0/word665 memory_8_0/word666 memory_8_0/word667 memory_8_0/word668 memory_8_0/word669
+ memory_8_0/word670 memory_8_0/word671 memory_8_0/word672 memory_8_0/word673 memory_8_0/word674
+ memory_8_0/word675 memory_8_0/word676 memory_8_0/word677 memory_8_0/word678 memory_8_0/word679
+ memory_8_0/word680 memory_8_0/word681 memory_8_0/word682 memory_8_0/word683 memory_8_0/word684
+ memory_8_0/word685 memory_8_0/word686 memory_8_0/word687 memory_8_0/word688 memory_8_0/word689
+ memory_8_0/word690 memory_8_0/word691 memory_8_0/word692 memory_8_0/word693 memory_8_0/word694
+ memory_8_0/word695 memory_8_0/word696 memory_8_0/word697 memory_8_0/word698 memory_8_0/word699
+ memory_8_0/word700 memory_8_0/word701 memory_8_0/word702 memory_8_0/word703 memory_8_0/word704
+ memory_8_0/word705 memory_8_0/word706 memory_8_0/word707 memory_8_0/word708 memory_8_0/word709
+ memory_8_0/word710 memory_8_0/word711 memory_8_0/word712 memory_8_0/word713 memory_8_0/word714
+ memory_8_0/word715 memory_8_0/word716 memory_8_0/word717 memory_8_0/word718 memory_8_0/word719
+ memory_8_0/word720 memory_8_0/word721 memory_8_0/word722 memory_8_0/word723 memory_8_0/word724
+ memory_8_0/word725 memory_8_0/word726 memory_8_0/word727 memory_8_0/word728 memory_8_0/word729
+ memory_8_0/word730 memory_8_0/word731 memory_8_0/word732 memory_8_0/word733 memory_8_0/word734
+ memory_8_0/word735 memory_8_0/word736 memory_8_0/word737 memory_8_0/word738 memory_8_0/word739
+ memory_8_0/word740 memory_8_0/word741 memory_8_0/word742 memory_8_0/word743 memory_8_0/word744
+ memory_8_0/word745 memory_8_0/word746 memory_8_0/word747 memory_8_0/word748 memory_8_0/word749
+ memory_8_0/word750 memory_8_0/word751 memory_8_0/word752 memory_8_0/word753 memory_8_0/word754
+ memory_8_0/word755 memory_8_0/word756 memory_8_0/word757 memory_8_0/word758 memory_8_0/word759
+ memory_8_0/word760 memory_8_0/word761 memory_8_0/word762 memory_8_0/word763 memory_8_0/word764
+ memory_8_0/word765 memory_8_0/word766 memory_8_0/word767 memory_8_0/word768 memory_8_0/word769
+ memory_8_0/word770 memory_8_0/word771 memory_8_0/word772 memory_8_0/word773 memory_8_0/word774
+ memory_8_0/word775 memory_8_0/word776 memory_8_0/word777 memory_8_0/word778 memory_8_0/word779
+ memory_8_0/word780 memory_8_0/word781 memory_8_0/word782 memory_8_0/word783 memory_8_0/word784
+ memory_8_0/word785 memory_8_0/word786 memory_8_0/word787 memory_8_0/word788 memory_8_0/word789
+ memory_8_0/word790 memory_8_0/word791 memory_8_0/word792 memory_8_0/word793 memory_8_0/word794
+ memory_8_0/word795 memory_8_0/word796 memory_8_0/word797 memory_8_0/word798 memory_8_0/word799
+ memory_8_0/word800 memory_8_0/word801 memory_8_0/word802 memory_8_0/word803 memory_8_0/word804
+ memory_8_0/word805 memory_8_0/word806 memory_8_0/word807 memory_8_0/word808 memory_8_0/word809
+ memory_8_0/word810 memory_8_0/word811 memory_8_0/word812 memory_8_0/word813 memory_8_0/word814
+ memory_8_0/word815 memory_8_0/word816 memory_8_0/word817 memory_8_0/word818 memory_8_0/word819
+ memory_8_0/word820 memory_8_0/word821 memory_8_0/word822 memory_8_0/word823 memory_8_0/word824
+ memory_8_0/word825 memory_8_0/word826 memory_8_0/word827 memory_8_0/word828 memory_8_0/word829
+ memory_8_0/word830 memory_8_0/word831 memory_8_0/word832 memory_8_0/word833 memory_8_0/word834
+ memory_8_0/word835 memory_8_0/word836 memory_8_0/word837 memory_8_0/word838 memory_8_0/word839
+ memory_8_0/word840 memory_8_0/word841 memory_8_0/word842 memory_8_0/word843 memory_8_0/word844
+ memory_8_0/word845 memory_8_0/word846 memory_8_0/word847 memory_8_0/word848 memory_8_0/word849
+ memory_8_0/word850 memory_8_0/word851 memory_8_0/word852 memory_8_0/word853 memory_8_0/word854
+ memory_8_0/word855 memory_8_0/word856 memory_8_0/word857 memory_8_0/word858 memory_8_0/word859
+ memory_8_0/word860 memory_8_0/word861 memory_8_0/word862 memory_8_0/word863 memory_8_0/word864
+ memory_8_0/word865 memory_8_0/word866 memory_8_0/word867 memory_8_0/word868 memory_8_0/word869
+ memory_8_0/word870 memory_8_0/word871 memory_8_0/word872 memory_8_0/word873 memory_8_0/word874
+ memory_8_0/word875 memory_8_0/word876 memory_8_0/word877 memory_8_0/word878 memory_8_0/word879
+ memory_8_0/word880 memory_8_0/word881 memory_8_0/word882 memory_8_0/word883 memory_8_0/word884
+ memory_8_0/word885 memory_8_0/word886 memory_8_0/word887 memory_8_0/word888 memory_8_0/word889
+ memory_8_0/word890 memory_8_0/word891 memory_8_0/word892 memory_8_0/word893 memory_8_0/word894
+ memory_8_0/word895 memory_8_0/word896 memory_8_0/word897 memory_8_0/word898 memory_8_0/word899
+ memory_8_0/word900 memory_8_0/word901 memory_8_0/word902 memory_8_0/word903 memory_8_0/word904
+ memory_8_0/word905 memory_8_0/word906 memory_8_0/word907 memory_8_0/word908 memory_8_0/word909
+ memory_8_0/word910 memory_8_0/word911 memory_8_0/word912 memory_8_0/word913 memory_8_0/word914
+ memory_8_0/word915 memory_8_0/word916 memory_8_0/word917 memory_8_0/word918 memory_8_0/word919
+ memory_8_0/word920 memory_8_0/word921 memory_8_0/word922 memory_8_0/word923 memory_8_0/word924
+ memory_8_0/word925 memory_8_0/word926 memory_8_0/word927 memory_8_0/word928 memory_8_0/word929
+ memory_8_0/word930 memory_8_0/word931 memory_8_0/word932 memory_8_0/word933 memory_8_0/word934
+ memory_8_0/word935 memory_8_0/word936 memory_8_0/word937 memory_8_0/word938 memory_8_0/word939
+ memory_8_0/word940 memory_8_0/word941 memory_8_0/word942 memory_8_0/word943 memory_8_0/word944
+ memory_8_0/word945 memory_8_0/word946 memory_8_0/word947 memory_8_0/word948 memory_8_0/word949
+ memory_8_0/word950 memory_8_0/word951 memory_8_0/word952 memory_8_0/word953 memory_8_0/word954
+ memory_8_0/word955 memory_8_0/word956 memory_8_0/word957 memory_8_0/word958 memory_8_0/word959
+ memory_8_0/word960 memory_8_0/word961 memory_8_0/word962 memory_8_0/word963 memory_8_0/word964
+ memory_8_0/word965 memory_8_0/word966 memory_8_0/word967 memory_8_0/word968 memory_8_0/word969
+ memory_8_0/word970 memory_8_0/word971 memory_8_0/word972 memory_8_0/word973 memory_8_0/word974
+ memory_8_0/word975 memory_8_0/word976 memory_8_0/word977 memory_8_0/word978 memory_8_0/word979
+ memory_8_0/word980 memory_8_0/word981 memory_8_0/word982 memory_8_0/word983 memory_8_0/word984
+ memory_8_0/word985 memory_8_0/word986 memory_8_0/word987 memory_8_0/word988 memory_8_0/word989
+ memory_8_0/word990 memory_8_0/word991 memory_8_0/word992 memory_8_0/word993 memory_8_0/word994
+ memory_8_0/word995 memory_8_0/word996 memory_8_0/word997 memory_8_0/word998 memory_8_0/word999
+ memory_8_0/word1000 memory_8_0/word1001 memory_8_0/word1002 memory_8_0/word1003
+ memory_8_0/word1004 memory_8_0/word1005 memory_8_0/word1006 memory_8_0/word1007
+ memory_8_0/word1008 memory_8_0/word1009 memory_8_0/word1010 memory_8_0/word1011
+ memory_8_0/word1012 memory_8_0/word1013 memory_8_0/word1014 memory_8_0/word1015
+ memory_8_0/word1016 memory_8_0/word1017 memory_8_0/word1018 memory_8_0/word1019
+ memory_8_0/word1020 memory_8_0/word1021 memory_8_0/word1022 memory_8_0/word1023
+ inv_6/A inv_7/A inv_3/A inv_2/A inv_5/A inv_4/A inv_9/A inv_8/A inv_9/GND inv_9/VDD
+ memory_8
Xmux4_0 mux4_0/I1 mux4_0/I2 mux4_0/I3 Freq0 inv_0/Y Freq1 inv_1/Y mux4_0/Y inv_9/VDD
+ mux4_0/I0 inv_9/GND mux4
Xinv_0 inv_9/VDD inv_9/GND Freq0 inv_0/Y inv
Xinv_1 inv_9/VDD inv_9/GND Freq1 inv_1/Y inv
Xcounter_8_0 mux4_0/Y decoder_8_0/A0 decoder_8_0/A2 decoder_8_0/A3 decoder_8_0/A4
+ decoder_8_0/A5 decoder_8_0/A6 decoder_8_0/A7 inv_9/GND decoder_8_0/A1 inv_9/VDD
+ counter_8
Xinv_2 inv_9/VDD inv_9/GND inv_2/A Y4 inv
Xinv_3 inv_9/VDD inv_9/GND inv_3/A Y5 inv
Xdecoder_8_0 decoder_8_0/A0 decoder_8_0/A1 decoder_8_0/A2 decoder_8_0/A3 decoder_8_0/A4
+ decoder_8_0/A5 decoder_8_0/A6 memory_8_0/word0 memory_8_0/word1 memory_8_0/word2
+ memory_8_0/word3 memory_8_0/word4 memory_8_0/word5 memory_8_0/word6 memory_8_0/word7
+ memory_8_0/word8 memory_8_0/word9 memory_8_0/word10 memory_8_0/word11 memory_8_0/word12
+ memory_8_0/word13 memory_8_0/word14 memory_8_0/word15 memory_8_0/word16 memory_8_0/word17
+ memory_8_0/word18 memory_8_0/word19 memory_8_0/word20 memory_8_0/word21 memory_8_0/word22
+ memory_8_0/word23 memory_8_0/word24 memory_8_0/word25 memory_8_0/word26 memory_8_0/word27
+ memory_8_0/word28 memory_8_0/word29 memory_8_0/word30 memory_8_0/word31 memory_8_0/word32
+ memory_8_0/word33 memory_8_0/word34 memory_8_0/word35 memory_8_0/word36 memory_8_0/word37
+ memory_8_0/word38 memory_8_0/word39 memory_8_0/word40 memory_8_0/word41 memory_8_0/word42
+ memory_8_0/word43 memory_8_0/word44 memory_8_0/word45 memory_8_0/word46 memory_8_0/word47
+ memory_8_0/word48 memory_8_0/word49 memory_8_0/word50 memory_8_0/word51 memory_8_0/word52
+ memory_8_0/word53 memory_8_0/word54 memory_8_0/word55 memory_8_0/word56 memory_8_0/word57
+ memory_8_0/word58 memory_8_0/word59 memory_8_0/word60 memory_8_0/word61 memory_8_0/word62
+ memory_8_0/word63 memory_8_0/word64 memory_8_0/word65 memory_8_0/word66 memory_8_0/word67
+ memory_8_0/word68 memory_8_0/word69 memory_8_0/word70 memory_8_0/word71 memory_8_0/word72
+ memory_8_0/word73 memory_8_0/word74 memory_8_0/word75 memory_8_0/word76 memory_8_0/word77
+ memory_8_0/word78 memory_8_0/word79 memory_8_0/word80 memory_8_0/word81 memory_8_0/word82
+ memory_8_0/word83 memory_8_0/word84 memory_8_0/word85 memory_8_0/word86 memory_8_0/word87
+ memory_8_0/word88 memory_8_0/word89 memory_8_0/word90 memory_8_0/word91 memory_8_0/word92
+ memory_8_0/word93 memory_8_0/word94 memory_8_0/word95 memory_8_0/word96 memory_8_0/word97
+ memory_8_0/word98 memory_8_0/word99 memory_8_0/word100 memory_8_0/word101 memory_8_0/word102
+ memory_8_0/word103 memory_8_0/word104 memory_8_0/word105 memory_8_0/word106 memory_8_0/word107
+ memory_8_0/word108 memory_8_0/word109 memory_8_0/word110 memory_8_0/word111 memory_8_0/word112
+ memory_8_0/word113 memory_8_0/word114 memory_8_0/word115 memory_8_0/word116 memory_8_0/word117
+ memory_8_0/word118 memory_8_0/word119 memory_8_0/word120 memory_8_0/word121 memory_8_0/word122
+ memory_8_0/word123 memory_8_0/word124 memory_8_0/word125 memory_8_0/word126 memory_8_0/word127
+ memory_8_0/word128 memory_8_0/word129 memory_8_0/word130 memory_8_0/word131 memory_8_0/word132
+ memory_8_0/word133 memory_8_0/word134 memory_8_0/word135 memory_8_0/word136 memory_8_0/word137
+ memory_8_0/word138 memory_8_0/word139 memory_8_0/word140 memory_8_0/word141 memory_8_0/word142
+ memory_8_0/word143 memory_8_0/word144 memory_8_0/word145 memory_8_0/word146 memory_8_0/word147
+ memory_8_0/word148 memory_8_0/word149 memory_8_0/word150 memory_8_0/word151 memory_8_0/word152
+ memory_8_0/word153 memory_8_0/word154 memory_8_0/word155 memory_8_0/word156 memory_8_0/word157
+ memory_8_0/word158 memory_8_0/word159 memory_8_0/word160 memory_8_0/word161 memory_8_0/word162
+ memory_8_0/word163 memory_8_0/word164 memory_8_0/word165 memory_8_0/word166 memory_8_0/word167
+ memory_8_0/word168 memory_8_0/word169 memory_8_0/word170 memory_8_0/word171 memory_8_0/word172
+ memory_8_0/word173 memory_8_0/word174 memory_8_0/word175 memory_8_0/word176 memory_8_0/word177
+ memory_8_0/word178 memory_8_0/word179 memory_8_0/word180 memory_8_0/word181 memory_8_0/word182
+ memory_8_0/word183 memory_8_0/word184 memory_8_0/word185 memory_8_0/word186 memory_8_0/word187
+ memory_8_0/word188 memory_8_0/word189 memory_8_0/word190 memory_8_0/word191 memory_8_0/word192
+ memory_8_0/word193 memory_8_0/word194 memory_8_0/word195 memory_8_0/word196 memory_8_0/word197
+ memory_8_0/word198 memory_8_0/word199 memory_8_0/word200 memory_8_0/word201 memory_8_0/word202
+ memory_8_0/word203 memory_8_0/word204 memory_8_0/word205 memory_8_0/word206 memory_8_0/word207
+ memory_8_0/word208 memory_8_0/word209 memory_8_0/word210 memory_8_0/word211 memory_8_0/word212
+ memory_8_0/word213 memory_8_0/word214 memory_8_0/word215 memory_8_0/word216 memory_8_0/word217
+ memory_8_0/word218 memory_8_0/word219 memory_8_0/word220 memory_8_0/word221 memory_8_0/word222
+ memory_8_0/word223 memory_8_0/word224 memory_8_0/word225 memory_8_0/word226 memory_8_0/word227
+ memory_8_0/word228 memory_8_0/word229 memory_8_0/word230 memory_8_0/word231 memory_8_0/word232
+ memory_8_0/word233 memory_8_0/word234 memory_8_0/word235 memory_8_0/word236 memory_8_0/word237
+ memory_8_0/word238 memory_8_0/word239 memory_8_0/word240 memory_8_0/word241 memory_8_0/word242
+ memory_8_0/word243 memory_8_0/word244 memory_8_0/word245 memory_8_0/word246 memory_8_0/word247
+ memory_8_0/word248 memory_8_0/word249 memory_8_0/word250 memory_8_0/word251 memory_8_0/word252
+ memory_8_0/word253 memory_8_0/word254 memory_8_0/word255 memory_8_0/word256 memory_8_0/word257
+ memory_8_0/word258 memory_8_0/word259 memory_8_0/word260 memory_8_0/word261 memory_8_0/word262
+ memory_8_0/word263 memory_8_0/word264 memory_8_0/word265 memory_8_0/word266 memory_8_0/word267
+ memory_8_0/word268 memory_8_0/word269 memory_8_0/word270 memory_8_0/word271 memory_8_0/word272
+ memory_8_0/word273 memory_8_0/word274 memory_8_0/word275 memory_8_0/word276 memory_8_0/word277
+ memory_8_0/word278 memory_8_0/word279 memory_8_0/word280 memory_8_0/word281 memory_8_0/word282
+ memory_8_0/word283 memory_8_0/word284 memory_8_0/word285 memory_8_0/word286 memory_8_0/word287
+ memory_8_0/word288 memory_8_0/word289 memory_8_0/word290 memory_8_0/word291 memory_8_0/word292
+ memory_8_0/word293 memory_8_0/word294 memory_8_0/word295 memory_8_0/word296 memory_8_0/word297
+ memory_8_0/word298 memory_8_0/word299 memory_8_0/word300 memory_8_0/word301 memory_8_0/word302
+ memory_8_0/word303 memory_8_0/word304 memory_8_0/word305 memory_8_0/word306 memory_8_0/word307
+ memory_8_0/word308 memory_8_0/word309 memory_8_0/word310 memory_8_0/word311 memory_8_0/word312
+ memory_8_0/word313 memory_8_0/word314 memory_8_0/word315 memory_8_0/word316 memory_8_0/word317
+ memory_8_0/word318 memory_8_0/word319 memory_8_0/word320 memory_8_0/word321 memory_8_0/word322
+ memory_8_0/word323 memory_8_0/word324 memory_8_0/word325 memory_8_0/word326 memory_8_0/word327
+ memory_8_0/word328 memory_8_0/word329 memory_8_0/word330 memory_8_0/word331 memory_8_0/word332
+ memory_8_0/word333 memory_8_0/word334 memory_8_0/word335 memory_8_0/word336 memory_8_0/word337
+ memory_8_0/word338 memory_8_0/word339 memory_8_0/word340 memory_8_0/word341 memory_8_0/word342
+ memory_8_0/word343 memory_8_0/word344 memory_8_0/word345 memory_8_0/word346 memory_8_0/word347
+ memory_8_0/word348 memory_8_0/word349 memory_8_0/word350 memory_8_0/word351 memory_8_0/word352
+ memory_8_0/word353 memory_8_0/word354 memory_8_0/word355 memory_8_0/word356 memory_8_0/word357
+ memory_8_0/word358 memory_8_0/word359 memory_8_0/word360 memory_8_0/word361 memory_8_0/word362
+ memory_8_0/word363 memory_8_0/word364 memory_8_0/word365 memory_8_0/word366 memory_8_0/word367
+ memory_8_0/word368 memory_8_0/word369 memory_8_0/word370 memory_8_0/word371 memory_8_0/word372
+ memory_8_0/word373 memory_8_0/word374 memory_8_0/word375 memory_8_0/word376 memory_8_0/word377
+ memory_8_0/word378 memory_8_0/word379 memory_8_0/word380 memory_8_0/word381 memory_8_0/word382
+ memory_8_0/word383 memory_8_0/word384 memory_8_0/word385 memory_8_0/word386 memory_8_0/word387
+ memory_8_0/word388 memory_8_0/word389 memory_8_0/word390 memory_8_0/word391 memory_8_0/word392
+ memory_8_0/word393 memory_8_0/word394 memory_8_0/word395 memory_8_0/word396 memory_8_0/word397
+ memory_8_0/word398 memory_8_0/word399 memory_8_0/word400 memory_8_0/word401 memory_8_0/word402
+ memory_8_0/word403 memory_8_0/word404 memory_8_0/word405 memory_8_0/word406 memory_8_0/word407
+ memory_8_0/word408 memory_8_0/word409 memory_8_0/word410 memory_8_0/word411 memory_8_0/word412
+ memory_8_0/word413 memory_8_0/word414 memory_8_0/word415 memory_8_0/word416 memory_8_0/word417
+ memory_8_0/word418 memory_8_0/word419 memory_8_0/word420 memory_8_0/word421 memory_8_0/word422
+ memory_8_0/word423 memory_8_0/word424 memory_8_0/word425 memory_8_0/word426 memory_8_0/word427
+ memory_8_0/word428 memory_8_0/word429 memory_8_0/word430 memory_8_0/word431 memory_8_0/word432
+ memory_8_0/word433 memory_8_0/word434 memory_8_0/word435 memory_8_0/word436 memory_8_0/word437
+ memory_8_0/word438 memory_8_0/word439 memory_8_0/word440 memory_8_0/word441 memory_8_0/word442
+ memory_8_0/word443 memory_8_0/word444 memory_8_0/word445 memory_8_0/word446 memory_8_0/word447
+ memory_8_0/word448 memory_8_0/word449 memory_8_0/word450 memory_8_0/word451 memory_8_0/word452
+ memory_8_0/word453 memory_8_0/word454 memory_8_0/word455 memory_8_0/word456 memory_8_0/word457
+ memory_8_0/word458 memory_8_0/word459 memory_8_0/word460 memory_8_0/word461 memory_8_0/word462
+ memory_8_0/word463 memory_8_0/word464 memory_8_0/word465 memory_8_0/word466 memory_8_0/word467
+ memory_8_0/word468 memory_8_0/word469 memory_8_0/word470 memory_8_0/word471 memory_8_0/word472
+ memory_8_0/word473 memory_8_0/word474 memory_8_0/word475 memory_8_0/word476 memory_8_0/word477
+ memory_8_0/word478 memory_8_0/word479 memory_8_0/word480 memory_8_0/word481 memory_8_0/word482
+ memory_8_0/word483 memory_8_0/word484 memory_8_0/word485 memory_8_0/word486 memory_8_0/word487
+ memory_8_0/word488 memory_8_0/word489 memory_8_0/word490 memory_8_0/word491 memory_8_0/word492
+ memory_8_0/word493 memory_8_0/word494 memory_8_0/word495 memory_8_0/word496 memory_8_0/word497
+ memory_8_0/word498 memory_8_0/word499 memory_8_0/word500 memory_8_0/word501 memory_8_0/word502
+ memory_8_0/word503 memory_8_0/word504 memory_8_0/word505 memory_8_0/word506 memory_8_0/word507
+ memory_8_0/word508 memory_8_0/word509 memory_8_0/word510 memory_8_0/word511 memory_8_0/word512
+ memory_8_0/word513 memory_8_0/word514 memory_8_0/word515 memory_8_0/word516 memory_8_0/word517
+ memory_8_0/word518 memory_8_0/word519 memory_8_0/word520 memory_8_0/word521 memory_8_0/word522
+ memory_8_0/word523 memory_8_0/word524 memory_8_0/word525 memory_8_0/word526 memory_8_0/word527
+ memory_8_0/word528 memory_8_0/word529 memory_8_0/word530 memory_8_0/word531 memory_8_0/word532
+ memory_8_0/word533 memory_8_0/word534 memory_8_0/word535 memory_8_0/word536 memory_8_0/word537
+ memory_8_0/word538 memory_8_0/word539 memory_8_0/word540 memory_8_0/word541 memory_8_0/word542
+ memory_8_0/word543 memory_8_0/word544 memory_8_0/word545 memory_8_0/word546 memory_8_0/word547
+ memory_8_0/word548 memory_8_0/word549 memory_8_0/word550 memory_8_0/word551 memory_8_0/word552
+ memory_8_0/word553 memory_8_0/word554 memory_8_0/word555 memory_8_0/word556 memory_8_0/word557
+ memory_8_0/word558 memory_8_0/word559 memory_8_0/word560 memory_8_0/word561 memory_8_0/word562
+ memory_8_0/word563 memory_8_0/word564 memory_8_0/word565 memory_8_0/word566 memory_8_0/word567
+ memory_8_0/word568 memory_8_0/word569 memory_8_0/word570 memory_8_0/word571 memory_8_0/word572
+ memory_8_0/word573 memory_8_0/word574 memory_8_0/word575 memory_8_0/word576 memory_8_0/word577
+ memory_8_0/word578 memory_8_0/word579 memory_8_0/word580 memory_8_0/word581 memory_8_0/word582
+ memory_8_0/word583 memory_8_0/word584 memory_8_0/word585 memory_8_0/word586 memory_8_0/word587
+ memory_8_0/word588 memory_8_0/word589 memory_8_0/word590 memory_8_0/word591 memory_8_0/word592
+ memory_8_0/word593 memory_8_0/word594 memory_8_0/word595 memory_8_0/word596 memory_8_0/word597
+ memory_8_0/word598 memory_8_0/word599 memory_8_0/word600 memory_8_0/word601 memory_8_0/word602
+ memory_8_0/word603 memory_8_0/word604 memory_8_0/word605 memory_8_0/word606 memory_8_0/word607
+ memory_8_0/word608 memory_8_0/word609 memory_8_0/word610 memory_8_0/word611 memory_8_0/word612
+ memory_8_0/word613 memory_8_0/word614 memory_8_0/word615 memory_8_0/word616 memory_8_0/word617
+ memory_8_0/word618 memory_8_0/word619 memory_8_0/word620 memory_8_0/word621 memory_8_0/word622
+ memory_8_0/word623 memory_8_0/word624 memory_8_0/word625 memory_8_0/word626 memory_8_0/word627
+ memory_8_0/word628 memory_8_0/word629 memory_8_0/word630 memory_8_0/word631 memory_8_0/word632
+ memory_8_0/word633 memory_8_0/word634 memory_8_0/word635 memory_8_0/word636 memory_8_0/word637
+ memory_8_0/word638 memory_8_0/word639 memory_8_0/word640 memory_8_0/word641 memory_8_0/word642
+ memory_8_0/word643 memory_8_0/word644 memory_8_0/word645 memory_8_0/word646 memory_8_0/word647
+ memory_8_0/word648 memory_8_0/word649 memory_8_0/word650 memory_8_0/word651 memory_8_0/word652
+ memory_8_0/word653 memory_8_0/word654 memory_8_0/word655 memory_8_0/word656 memory_8_0/word657
+ memory_8_0/word658 memory_8_0/word659 memory_8_0/word660 memory_8_0/word661 memory_8_0/word662
+ memory_8_0/word663 memory_8_0/word664 memory_8_0/word665 memory_8_0/word666 memory_8_0/word667
+ memory_8_0/word668 memory_8_0/word669 memory_8_0/word670 memory_8_0/word671 memory_8_0/word672
+ memory_8_0/word673 memory_8_0/word674 memory_8_0/word675 memory_8_0/word676 memory_8_0/word677
+ memory_8_0/word678 memory_8_0/word679 memory_8_0/word680 memory_8_0/word681 memory_8_0/word682
+ memory_8_0/word683 memory_8_0/word684 memory_8_0/word685 memory_8_0/word686 memory_8_0/word687
+ memory_8_0/word688 memory_8_0/word689 memory_8_0/word690 memory_8_0/word691 memory_8_0/word692
+ memory_8_0/word693 memory_8_0/word694 memory_8_0/word695 memory_8_0/word696 memory_8_0/word697
+ memory_8_0/word698 memory_8_0/word699 memory_8_0/word700 memory_8_0/word701 memory_8_0/word702
+ memory_8_0/word703 memory_8_0/word704 memory_8_0/word705 memory_8_0/word706 memory_8_0/word707
+ memory_8_0/word708 memory_8_0/word709 memory_8_0/word710 memory_8_0/word711 memory_8_0/word712
+ memory_8_0/word713 memory_8_0/word714 memory_8_0/word715 memory_8_0/word716 memory_8_0/word717
+ memory_8_0/word718 memory_8_0/word719 memory_8_0/word720 memory_8_0/word721 memory_8_0/word722
+ memory_8_0/word723 memory_8_0/word724 memory_8_0/word725 memory_8_0/word726 memory_8_0/word727
+ memory_8_0/word728 memory_8_0/word729 memory_8_0/word730 memory_8_0/word731 memory_8_0/word732
+ memory_8_0/word733 memory_8_0/word734 memory_8_0/word735 memory_8_0/word736 memory_8_0/word737
+ memory_8_0/word738 memory_8_0/word739 memory_8_0/word740 memory_8_0/word741 memory_8_0/word742
+ memory_8_0/word743 memory_8_0/word744 memory_8_0/word745 memory_8_0/word746 memory_8_0/word747
+ memory_8_0/word748 memory_8_0/word749 memory_8_0/word750 memory_8_0/word751 memory_8_0/word752
+ memory_8_0/word753 memory_8_0/word754 memory_8_0/word755 memory_8_0/word756 memory_8_0/word757
+ memory_8_0/word758 memory_8_0/word759 memory_8_0/word760 memory_8_0/word761 memory_8_0/word762
+ memory_8_0/word763 memory_8_0/word764 memory_8_0/word765 memory_8_0/word766 memory_8_0/word767
+ memory_8_0/word768 memory_8_0/word769 memory_8_0/word770 memory_8_0/word771 memory_8_0/word772
+ memory_8_0/word773 memory_8_0/word774 memory_8_0/word775 memory_8_0/word776 memory_8_0/word777
+ memory_8_0/word778 memory_8_0/word779 memory_8_0/word780 memory_8_0/word781 memory_8_0/word782
+ memory_8_0/word783 memory_8_0/word784 memory_8_0/word785 memory_8_0/word786 memory_8_0/word787
+ memory_8_0/word788 memory_8_0/word789 memory_8_0/word790 memory_8_0/word791 memory_8_0/word792
+ memory_8_0/word793 memory_8_0/word794 memory_8_0/word795 memory_8_0/word796 memory_8_0/word797
+ memory_8_0/word798 memory_8_0/word799 memory_8_0/word800 memory_8_0/word801 memory_8_0/word802
+ memory_8_0/word803 memory_8_0/word804 memory_8_0/word805 memory_8_0/word806 memory_8_0/word807
+ memory_8_0/word808 memory_8_0/word809 memory_8_0/word810 memory_8_0/word811 memory_8_0/word812
+ memory_8_0/word813 memory_8_0/word814 memory_8_0/word815 memory_8_0/word816 memory_8_0/word817
+ memory_8_0/word818 memory_8_0/word819 memory_8_0/word820 memory_8_0/word821 memory_8_0/word822
+ memory_8_0/word823 memory_8_0/word824 memory_8_0/word825 memory_8_0/word826 memory_8_0/word827
+ memory_8_0/word828 memory_8_0/word829 memory_8_0/word830 memory_8_0/word831 memory_8_0/word832
+ memory_8_0/word833 memory_8_0/word834 memory_8_0/word835 memory_8_0/word836 memory_8_0/word837
+ memory_8_0/word838 memory_8_0/word839 memory_8_0/word840 memory_8_0/word841 memory_8_0/word842
+ memory_8_0/word843 memory_8_0/word844 memory_8_0/word845 memory_8_0/word846 memory_8_0/word847
+ memory_8_0/word848 memory_8_0/word849 memory_8_0/word850 memory_8_0/word851 memory_8_0/word852
+ memory_8_0/word853 memory_8_0/word854 memory_8_0/word855 memory_8_0/word856 memory_8_0/word857
+ memory_8_0/word858 memory_8_0/word859 memory_8_0/word860 memory_8_0/word861 memory_8_0/word862
+ memory_8_0/word863 memory_8_0/word864 memory_8_0/word865 memory_8_0/word866 memory_8_0/word867
+ memory_8_0/word868 memory_8_0/word869 memory_8_0/word870 memory_8_0/word871 memory_8_0/word872
+ memory_8_0/word873 memory_8_0/word874 memory_8_0/word875 memory_8_0/word876 memory_8_0/word877
+ memory_8_0/word878 memory_8_0/word879 memory_8_0/word880 memory_8_0/word881 memory_8_0/word882
+ memory_8_0/word883 memory_8_0/word884 memory_8_0/word885 memory_8_0/word886 memory_8_0/word887
+ memory_8_0/word888 memory_8_0/word889 memory_8_0/word890 memory_8_0/word891 memory_8_0/word892
+ memory_8_0/word893 memory_8_0/word894 memory_8_0/word895 memory_8_0/word896 memory_8_0/word897
+ memory_8_0/word898 memory_8_0/word899 memory_8_0/word900 memory_8_0/word901 memory_8_0/word902
+ memory_8_0/word903 memory_8_0/word904 memory_8_0/word905 memory_8_0/word906 memory_8_0/word907
+ memory_8_0/word908 memory_8_0/word909 memory_8_0/word910 memory_8_0/word911 memory_8_0/word912
+ memory_8_0/word913 memory_8_0/word914 memory_8_0/word915 memory_8_0/word916 memory_8_0/word917
+ memory_8_0/word918 memory_8_0/word919 memory_8_0/word920 memory_8_0/word921 memory_8_0/word922
+ memory_8_0/word923 memory_8_0/word924 memory_8_0/word925 memory_8_0/word926 memory_8_0/word927
+ memory_8_0/word928 memory_8_0/word929 memory_8_0/word930 memory_8_0/word931 memory_8_0/word932
+ memory_8_0/word933 memory_8_0/word934 memory_8_0/word935 memory_8_0/word936 memory_8_0/word937
+ memory_8_0/word938 memory_8_0/word939 memory_8_0/word940 memory_8_0/word941 memory_8_0/word942
+ memory_8_0/word943 memory_8_0/word944 memory_8_0/word945 memory_8_0/word946 memory_8_0/word947
+ memory_8_0/word948 memory_8_0/word949 memory_8_0/word950 memory_8_0/word951 memory_8_0/word952
+ memory_8_0/word953 memory_8_0/word954 memory_8_0/word955 memory_8_0/word956 memory_8_0/word957
+ memory_8_0/word958 memory_8_0/word959 memory_8_0/word960 memory_8_0/word961 memory_8_0/word962
+ memory_8_0/word963 memory_8_0/word964 memory_8_0/word965 memory_8_0/word966 memory_8_0/word967
+ memory_8_0/word968 memory_8_0/word969 memory_8_0/word970 memory_8_0/word971 memory_8_0/word972
+ memory_8_0/word973 memory_8_0/word974 memory_8_0/word975 memory_8_0/word976 memory_8_0/word977
+ memory_8_0/word978 memory_8_0/word979 memory_8_0/word980 memory_8_0/word981 memory_8_0/word982
+ memory_8_0/word983 memory_8_0/word984 memory_8_0/word985 memory_8_0/word986 memory_8_0/word987
+ memory_8_0/word988 memory_8_0/word989 memory_8_0/word990 memory_8_0/word991 memory_8_0/word992
+ memory_8_0/word993 memory_8_0/word994 memory_8_0/word995 memory_8_0/word996 memory_8_0/word997
+ memory_8_0/word998 memory_8_0/word999 memory_8_0/word1000 memory_8_0/word1001 memory_8_0/word1002
+ memory_8_0/word1003 memory_8_0/word1004 memory_8_0/word1005 memory_8_0/word1006
+ memory_8_0/word1007 memory_8_0/word1008 memory_8_0/word1009 memory_8_0/word1010
+ memory_8_0/word1011 memory_8_0/word1012 memory_8_0/word1013 memory_8_0/word1014
+ memory_8_0/word1015 memory_8_0/word1016 memory_8_0/word1017 memory_8_0/word1018
+ memory_8_0/word1019 memory_8_0/word1020 memory_8_0/word1021 memory_8_0/word1022
+ memory_8_0/word1023 inv_9/VDD inv_9/GND decoder_8_0/A7 Wave0 Wave1 decoder_8
Xinv_4 inv_9/VDD inv_9/GND inv_4/A Y2 inv
Xinv_5 inv_9/VDD inv_9/GND inv_5/A Y3 inv
Xinv_7 inv_9/VDD inv_9/GND inv_7/A Y6 inv
Xinv_6 inv_9/VDD inv_9/GND inv_6/A Y7 inv
Xcounter_4_0 CLK mux4_0/I0 mux4_0/I1 mux4_0/I2 mux4_0/I3 inv_9/GND inv_9/VDD counter_4
Xinv_8 inv_9/VDD inv_9/GND inv_8/A Y0 inv
Xinv_9 inv_9/VDD inv_9/GND inv_9/A Y1 inv
*.ends

