magic
tech sky130A
timestamp 1741623493
<< nwell >>
rect -2 197 323 488
<< nmos >>
rect 72 113 87 163
rect 126 113 141 163
rect 180 113 195 163
rect 234 113 249 163
<< pmos >>
rect 72 315 87 415
rect 126 315 141 415
rect 180 315 195 415
rect 234 315 249 415
<< ndiff >>
rect 36 155 72 163
rect 36 121 44 155
rect 61 121 72 155
rect 36 113 72 121
rect 87 155 126 163
rect 87 121 98 155
rect 115 121 126 155
rect 87 113 126 121
rect 141 155 180 163
rect 141 121 152 155
rect 169 121 180 155
rect 141 113 180 121
rect 195 155 234 163
rect 195 121 206 155
rect 223 121 234 155
rect 195 113 234 121
rect 249 155 285 163
rect 249 121 260 155
rect 277 121 285 155
rect 249 113 285 121
<< pdiff >>
rect 36 407 72 415
rect 36 323 44 407
rect 61 323 72 407
rect 36 315 72 323
rect 87 315 126 415
rect 141 407 180 415
rect 141 323 152 407
rect 169 323 180 407
rect 141 315 180 323
rect 195 315 234 415
rect 249 407 285 415
rect 249 323 260 407
rect 277 323 285 407
rect 249 315 285 323
<< ndiffc >>
rect 44 121 61 155
rect 98 121 115 155
rect 152 121 169 155
rect 206 121 223 155
rect 260 121 277 155
<< pdiffc >>
rect 44 323 61 407
rect 152 323 169 407
rect 260 323 277 407
<< psubdiff >>
rect 0 10 12 38
rect 309 10 321 38
<< nsubdiff >>
rect 16 442 28 470
rect 293 442 305 470
<< psubdiffcont >>
rect 12 10 309 38
<< nsubdiffcont >>
rect 28 442 293 470
<< poly >>
rect 72 415 87 428
rect 126 415 141 428
rect 180 415 195 428
rect 234 415 249 428
rect 72 290 87 315
rect 54 282 87 290
rect 54 265 62 282
rect 79 265 87 282
rect 54 257 87 265
rect 72 163 87 257
rect 126 250 141 315
rect 180 250 195 315
rect 108 242 141 250
rect 108 225 116 242
rect 133 225 141 242
rect 108 217 141 225
rect 162 242 195 250
rect 162 225 170 242
rect 187 225 195 242
rect 162 217 195 225
rect 126 163 141 217
rect 180 163 195 217
rect 234 298 249 315
rect 234 290 282 298
rect 234 273 257 290
rect 274 273 282 290
rect 234 265 282 273
rect 234 163 249 265
rect 72 100 87 113
rect 126 100 141 113
rect 180 100 195 113
rect 234 100 249 113
<< polycont >>
rect 62 265 79 282
rect 116 225 133 242
rect 170 225 187 242
rect 257 273 274 290
<< locali >>
rect 0 470 321 480
rect 0 442 28 470
rect 293 442 321 470
rect 0 432 321 442
rect 36 407 69 432
rect 36 323 44 407
rect 61 323 69 407
rect 36 315 69 323
rect 144 407 177 415
rect 144 323 152 407
rect 169 323 177 407
rect 54 282 87 290
rect 54 265 62 282
rect 79 265 87 282
rect 144 288 177 323
rect 252 407 285 432
rect 252 323 260 407
rect 277 323 285 407
rect 252 315 285 323
rect 249 290 282 298
rect 144 271 231 288
rect 54 257 87 265
rect 108 242 141 250
rect 108 225 116 242
rect 133 225 141 242
rect 108 217 141 225
rect 162 242 195 250
rect 162 225 170 242
rect 187 225 195 242
rect 162 217 195 225
rect 212 228 231 271
rect 249 273 257 290
rect 274 273 282 290
rect 249 265 282 273
rect 284 228 317 239
rect 212 206 317 228
rect 36 180 177 200
rect 36 155 69 180
rect 36 121 44 155
rect 61 121 69 155
rect 36 113 69 121
rect 90 155 123 163
rect 90 121 98 155
rect 115 121 123 155
rect 90 48 123 121
rect 144 155 177 180
rect 212 168 231 206
rect 144 121 152 155
rect 169 121 177 155
rect 144 84 177 121
rect 198 155 231 168
rect 198 121 206 155
rect 223 121 231 155
rect 198 113 231 121
rect 252 155 285 163
rect 252 121 260 155
rect 277 121 285 155
rect 252 84 285 121
rect 144 67 285 84
rect 0 38 321 48
rect 0 10 12 38
rect 309 10 321 38
rect 0 0 321 10
<< labels >>
flabel pdiff 72 365 72 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 195 365 195 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 249 365 249 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 126 363 126 363 1 FreeSerif 8 0 0 0 S$
flabel ndiff 87 135 87 135 1 FreeSerif 8 0 0 0 S$
flabel ndiff 126 137 126 137 1 FreeSerif 8 0 0 0 S$
flabel ndiff 180 137 180 137 1 FreeSerif 8 0 0 0 S$
flabel ndiff 249 138 249 138 1 FreeSerif 8 0 0 0 S$
flabel locali 249 265 282 298 0 FreeSerif 80 0 0 0 I1
port 1 nsew
flabel locali 162 217 195 250 0 FreeSerif 80 0 0 0 ~S0
port 14 nsew
flabel locali 108 217 141 250 0 FreeSerif 80 0 0 0 S0
port 4 nsew
flabel locali 54 257 87 290 0 FreeSerif 80 0 0 0 I0
port 2 nsew
flabel locali 284 206 317 239 0 FreeSerif 80 0 0 0 Y
port 11 nsew
flabel locali 0 432 321 480 0 FreeSerif 80 0 0 0 VDD!
port 9 nsew
flabel locali 0 0 321 48 0 FreeSerif 80 0 0 0 GND!
port 10 nsew
<< end >>
