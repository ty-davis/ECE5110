magic
tech sky130A
timestamp 1744679307
<< poly >>
rect -51 -17 792 0
rect -51 -88 792 -71
rect -51 -159 792 -142
rect -51 -230 792 -213
rect -51 -301 792 -284
rect -51 -372 792 -355
rect -51 -443 792 -426
rect -51 -514 792 -497
rect -51 -585 792 -568
rect -51 -656 792 -639
rect -51 -727 792 -710
rect -51 -798 792 -781
rect -51 -869 792 -852
rect -51 -940 792 -923
rect -51 -1011 792 -994
rect -51 -1082 792 -1065
rect -51 -1153 792 -1136
rect -51 -1224 792 -1207
rect -51 -1295 792 -1278
rect -51 -1366 792 -1349
rect -51 -1437 792 -1420
rect -51 -1508 792 -1491
rect -51 -1579 792 -1562
rect -51 -1650 792 -1633
rect -51 -1721 792 -1704
rect -51 -1792 792 -1775
rect -51 -1863 792 -1846
rect -51 -1934 792 -1917
rect -51 -2005 792 -1988
rect -51 -2076 792 -2059
rect -51 -2147 792 -2130
rect -51 -2218 792 -2201
rect -51 -2289 792 -2272
rect -51 -2360 792 -2343
rect -51 -2431 792 -2414
rect -51 -2502 792 -2485
rect -51 -2573 792 -2556
rect -51 -2644 792 -2627
rect -51 -2715 792 -2698
rect -51 -2786 792 -2769
rect -51 -2857 792 -2840
rect -51 -2928 792 -2911
rect -51 -2999 792 -2982
rect -51 -3070 792 -3053
rect -51 -3141 792 -3124
rect -51 -3212 792 -3195
rect -51 -3283 792 -3266
rect -51 -3354 792 -3337
rect -51 -3425 792 -3408
rect -51 -3496 792 -3479
rect -51 -3567 792 -3550
rect -51 -3638 792 -3621
rect -51 -3709 792 -3692
rect -51 -3780 792 -3763
rect -51 -3851 792 -3834
rect -51 -3922 792 -3905
rect -51 -3993 792 -3976
rect -51 -4064 792 -4047
rect -51 -4135 792 -4118
rect -51 -4206 792 -4189
rect -51 -4277 792 -4260
rect -51 -4348 792 -4331
rect -51 -4419 792 -4402
rect -51 -4490 792 -4473
rect -51 -4561 792 -4544
rect -51 -4632 792 -4615
rect -51 -4703 792 -4686
rect -51 -4774 792 -4757
rect -51 -4845 792 -4828
rect -51 -4916 792 -4899
rect -51 -4987 792 -4970
rect -51 -5058 792 -5041
rect -51 -5129 792 -5112
rect -51 -5200 792 -5183
rect -51 -5271 792 -5254
rect -51 -5342 792 -5325
rect -51 -5413 792 -5396
rect -51 -5484 792 -5467
rect -51 -5555 792 -5538
rect -51 -5626 792 -5609
rect -51 -5697 792 -5680
rect -51 -5768 792 -5751
rect -51 -5839 792 -5822
rect -51 -5910 792 -5893
rect -51 -5981 792 -5964
rect -51 -6052 792 -6035
rect -51 -6123 792 -6106
rect -51 -6194 792 -6177
rect -51 -6265 792 -6248
rect -51 -6336 792 -6319
rect -51 -6407 792 -6390
rect -51 -6478 792 -6461
rect -51 -6549 792 -6532
rect -51 -6620 792 -6603
rect -51 -6691 792 -6674
rect -51 -6762 792 -6745
rect -51 -6833 792 -6816
rect -51 -6904 792 -6887
rect -51 -6975 792 -6958
rect -51 -7046 792 -7029
rect -51 -7117 792 -7100
rect -51 -7188 792 -7171
rect -51 -7259 792 -7242
rect -51 -7330 792 -7313
rect -51 -7401 792 -7384
rect -51 -7472 792 -7455
rect -51 -7543 792 -7526
rect -51 -7614 792 -7597
rect -51 -7685 792 -7668
rect -51 -7756 792 -7739
rect -51 -7827 792 -7810
rect -51 -7898 792 -7881
rect -51 -7969 792 -7952
rect -51 -8040 792 -8023
rect -51 -8111 792 -8094
rect -51 -8182 792 -8165
rect -51 -8253 792 -8236
rect -51 -8324 792 -8307
rect -51 -8395 792 -8378
rect -51 -8466 792 -8449
rect -51 -8537 792 -8520
rect -51 -8608 792 -8591
rect -51 -8679 792 -8662
rect -51 -8750 792 -8733
rect -51 -8821 792 -8804
rect -51 -8892 792 -8875
rect -51 -8963 792 -8946
rect -51 -9034 792 -9017
<< locali >>
rect 0 -9088 33 41
rect 66 -9088 99 41
rect 132 -9088 165 41
rect 198 -9088 231 41
rect 264 -9088 297 41
rect 330 -9088 363 41
rect 396 -9088 429 41
rect 462 -9088 495 41
rect 528 -9088 561 41
rect 594 -9088 627 41
rect 660 -9088 693 41
rect 726 -9088 759 41
<< end >>