magic
tech sky130A
magscale 1 2
timestamp 1745496437
<< error_s >>
rect 60 145672 166 145682
<< nwell >>
rect -816 119516 -782 119552
rect 0 80 2914 118
<< locali >>
rect -114 146128 84 146176
rect -974 145854 -926 145860
rect -974 145818 -968 145854
rect -932 145818 -926 145854
rect -974 145626 -926 145818
rect -114 145628 -66 146128
rect 5758 146042 5814 146048
rect 5758 145998 5764 146042
rect 5808 145998 5814 146042
rect 36 145700 84 145818
rect 5758 145732 5814 145998
rect 6028 145992 6114 146048
rect 5660 145676 5814 145732
rect 5860 145626 6040 145706
rect -459 145434 -393 145567
rect -577 119909 -511 120090
rect -830 119563 -770 119564
rect -619 119563 -553 119782
rect -839 119552 -553 119563
rect -839 119516 -820 119552
rect -782 119516 -553 119552
rect -839 119504 -553 119516
rect 50 -84 106 140
rect 50 -128 56 -84
rect 100 -128 106 -84
rect 50 -134 106 -128
rect 5270 -924 5366 18
rect 5598 -134 5704 -78
rect 5828 -674 5894 -472
rect 6136 -674 6202 -472
rect 6444 -674 6510 -472
rect 6752 -564 6818 -362
rect 7060 -584 7126 -382
rect 7368 -592 7434 -390
rect 7676 -594 7742 -392
rect 7984 -598 8050 -396
rect 5270 -1020 5670 -924
<< viali >>
rect -968 145818 -932 145854
rect 5764 145998 5808 146042
rect 36 145818 84 145854
rect 5984 145992 6028 146048
rect -459 145567 -393 145621
rect -390 119936 -348 119976
rect -577 119855 -511 119909
rect -388 119628 -352 119670
rect -820 119516 -782 119552
rect -518 119462 -452 119528
rect -533 119223 -479 119277
rect -533 119115 -479 119169
rect -631 118767 -577 118821
rect -613 118365 -559 118419
rect -631 118131 -577 118185
rect -621 117735 -551 117805
rect -471 117316 -417 117370
rect 56 -128 100 -84
rect 6108 6 6174 60
rect 6440 9 6506 75
rect 6606 7 6672 73
rect 6938 13 7004 67
rect 7104 6 7170 60
rect 7436 6 7502 72
rect 7602 6 7668 60
rect 7934 9 8000 75
rect 5554 -134 5598 -78
rect 5733 -713 5787 -659
rect 6039 -715 6093 -661
rect 6341 -715 6395 -661
rect 6653 -713 6707 -659
rect 6967 -717 7021 -663
rect 7263 -723 7317 -669
rect 7565 -715 7619 -661
rect 7883 -715 7937 -661
<< metal1 >>
rect 5978 146048 6034 146060
rect 5752 146042 5984 146048
rect 5752 145998 5764 146042
rect 5808 145998 5984 146042
rect 5752 145992 5984 145998
rect 6028 145992 6034 146048
rect 5978 145980 6034 145992
rect -974 145860 -926 145866
rect -974 145854 96 145860
rect -974 145818 -968 145854
rect -932 145818 36 145854
rect 84 145818 96 145854
rect -974 145812 96 145818
rect -974 145806 -926 145812
rect -474 145627 -380 145634
rect -474 145561 -465 145627
rect -387 145561 -380 145627
rect -474 145554 -380 145561
rect -172 142385 -86 142396
rect -401 142319 -161 142385
rect -95 142319 -86 142385
rect -172 142310 -86 142319
rect -182 139130 -104 139138
rect -399 139064 -177 139130
rect -111 139064 -104 139130
rect -182 139058 -104 139064
rect -150 135919 -74 135932
rect -150 135917 -138 135919
rect -392 135868 -138 135917
rect -150 135867 -138 135868
rect -86 135867 -74 135919
rect -150 135856 -74 135867
rect -144 132659 -60 132668
rect -401 132593 -135 132659
rect -69 132593 -60 132659
rect -144 132582 -60 132593
rect -128 129425 -44 129434
rect -401 129359 -119 129425
rect -53 129359 -44 129425
rect -128 129350 -44 129359
rect -144 126183 -60 126192
rect -401 126117 -139 126183
rect -73 126117 -60 126183
rect -144 126108 -60 126117
rect -166 122951 -82 122960
rect -401 122885 -157 122951
rect -91 122885 -82 122951
rect -166 122876 -82 122885
rect -402 119976 -137 119988
rect -402 119936 -390 119976
rect -348 119936 -137 119976
rect -402 119922 -137 119936
rect -589 119909 -499 119915
rect -589 119855 -577 119909
rect -511 119873 -499 119909
rect -511 119855 -241 119873
rect -589 119849 -241 119855
rect -577 119807 -241 119849
rect -963 119670 -336 119680
rect -963 119628 -388 119670
rect -352 119628 -336 119670
rect -963 119614 -336 119628
rect -963 118549 -897 119614
rect -835 119552 -764 119569
rect -835 119516 -820 119552
rect -782 119516 -764 119552
rect -835 119498 -764 119516
rect -532 119534 -438 119540
rect -829 118656 -770 119498
rect -532 119456 -524 119534
rect -446 119456 -438 119534
rect -532 119450 -438 119456
rect -307 119283 -241 119807
rect -545 119277 -241 119283
rect -545 119223 -533 119277
rect -479 119223 -241 119277
rect -545 119217 -241 119223
rect -203 119175 -137 119922
rect -545 119169 -137 119175
rect -545 119115 -533 119169
rect -479 119115 -137 119169
rect -545 119109 -137 119115
rect -637 118827 -571 118833
rect -637 118755 -571 118761
rect -829 118597 -503 118656
rect -963 118483 -701 118549
rect -626 118425 -546 118432
rect -626 118359 -619 118425
rect -553 118359 -546 118425
rect -626 118352 -546 118359
rect -644 118191 -564 118198
rect -644 118125 -637 118191
rect -571 118125 -564 118191
rect -644 118118 -564 118125
rect -634 117811 -538 117818
rect -634 117729 -627 117811
rect -545 117729 -538 117811
rect -634 117722 -538 117729
rect -477 117376 -411 117382
rect -477 117304 -411 117310
rect -412 114390 -346 114400
rect -412 114316 -398 114390
rect -346 114316 -335 114365
rect -401 114299 -335 114316
rect -406 107894 -332 107904
rect -406 107814 -394 107894
rect -338 107814 -332 107894
rect -406 107802 -332 107814
rect 6088 80 6196 92
rect 6088 60 6198 80
rect 6088 6 6108 60
rect 6174 6 6198 60
rect 6088 -2 6198 6
rect 6428 75 6536 94
rect 6428 9 6440 75
rect 6506 9 6536 75
rect 6428 0 6536 9
rect 6592 73 6700 96
rect 6592 7 6606 73
rect 6672 7 6700 73
rect 6592 2 6700 7
rect 6920 67 7028 100
rect 6920 13 6938 67
rect 7004 13 7028 67
rect 6920 6 7028 13
rect 7090 66 7198 94
rect 7418 72 7526 92
rect 7090 60 7210 66
rect 7090 6 7104 60
rect 7170 6 7210 60
rect 6600 1 6678 2
rect 50 -78 106 -72
rect 5548 -78 5604 -66
rect 50 -84 5554 -78
rect 50 -128 56 -84
rect 100 -128 5554 -84
rect 50 -134 5554 -128
rect 5598 -134 5604 -78
rect 50 -140 106 -134
rect 5548 -146 5604 -134
rect 6108 -205 6174 -2
rect 5727 -271 6174 -205
rect 5727 -659 5793 -271
rect 6440 -311 6506 0
rect 5727 -713 5733 -659
rect 5787 -713 5793 -659
rect 5727 -725 5793 -713
rect 6033 -377 6506 -311
rect 6033 -661 6099 -377
rect 6606 -439 6672 1
rect 6033 -715 6039 -661
rect 6093 -715 6099 -661
rect 6033 -727 6099 -715
rect 6335 -505 6672 -439
rect 6335 -661 6401 -505
rect 6938 -523 7004 6
rect 7090 0 7210 6
rect 6829 -589 7004 -523
rect 7141 -466 7210 0
rect 7418 6 7436 72
rect 7502 6 7526 72
rect 7418 -2 7526 6
rect 7586 60 7694 94
rect 7930 81 8038 90
rect 7928 75 8038 81
rect 7586 6 7602 60
rect 7668 6 7694 60
rect 7586 0 7694 6
rect 7877 9 7934 75
rect 8000 9 8038 75
rect 6829 -653 6895 -589
rect 6335 -715 6341 -661
rect 6395 -715 6401 -661
rect 6335 -727 6401 -715
rect 6641 -659 6895 -653
rect 7141 -657 7207 -466
rect 6641 -713 6653 -659
rect 6707 -713 6895 -659
rect 6641 -719 6895 -713
rect 6955 -663 7207 -657
rect 7436 -663 7502 -2
rect 7602 -655 7668 0
rect 6955 -717 6967 -663
rect 7021 -717 7207 -663
rect 6955 -723 7207 -717
rect 7251 -669 7502 -663
rect 7251 -723 7263 -669
rect 7317 -723 7502 -669
rect 7553 -661 7668 -655
rect 7553 -715 7565 -661
rect 7619 -715 7668 -661
rect 7553 -721 7668 -715
rect 7877 -4 8038 9
rect 7877 -661 7943 -4
rect 7877 -715 7883 -661
rect 7937 -715 7943 -661
rect 7251 -729 7502 -723
rect 7877 -727 7943 -715
<< via1 >>
rect -465 145621 -387 145627
rect -465 145567 -459 145621
rect -459 145567 -393 145621
rect -393 145567 -387 145621
rect -465 145561 -387 145567
rect -161 142319 -95 142385
rect -177 139064 -111 139130
rect -138 135867 -86 135919
rect -135 132593 -69 132659
rect -119 129359 -53 129425
rect -139 126117 -73 126183
rect -157 122885 -91 122951
rect -524 119528 -446 119534
rect -524 119462 -518 119528
rect -518 119462 -452 119528
rect -452 119462 -446 119528
rect -524 119456 -446 119462
rect -637 118821 -571 118827
rect -637 118767 -631 118821
rect -631 118767 -577 118821
rect -577 118767 -571 118821
rect -637 118761 -571 118767
rect -619 118419 -553 118425
rect -619 118365 -613 118419
rect -613 118365 -559 118419
rect -559 118365 -553 118419
rect -619 118359 -553 118365
rect -637 118185 -571 118191
rect -637 118131 -631 118185
rect -631 118131 -577 118185
rect -577 118131 -571 118185
rect -637 118125 -571 118131
rect -627 117805 -545 117811
rect -627 117735 -621 117805
rect -621 117735 -551 117805
rect -551 117735 -545 117805
rect -627 117729 -545 117735
rect -477 117370 -411 117376
rect -477 117316 -471 117370
rect -471 117316 -417 117370
rect -417 117316 -411 117370
rect -477 117310 -411 117316
rect -398 114316 -346 114390
rect -401 111057 -335 111123
rect -394 107814 -338 107894
<< metal2 >>
rect 436 146748 502 146814
rect 700 146654 766 146720
rect 957 146626 1023 146635
rect 957 146560 1030 146626
rect -474 145627 -380 145634
rect -474 145561 -465 145627
rect -387 145561 -380 145627
rect 957 145622 1023 146560
rect 1222 146532 1289 146535
rect 1222 146466 1294 146532
rect 953 145566 962 145622
rect 1018 145566 1027 145622
rect 957 145561 1023 145566
rect -474 145554 -380 145561
rect -172 142385 -86 142396
rect -172 142319 -161 142385
rect -95 142319 -86 142385
rect 1222 142381 1289 146466
rect 1479 146436 1550 146442
rect 1479 146370 1562 146436
rect 1216 142324 1225 142381
rect 1286 142324 1295 142381
rect 1222 142319 1289 142324
rect -172 142310 -86 142319
rect -182 139130 -104 139138
rect -182 139064 -177 139130
rect -111 139064 -104 139130
rect -182 139058 -104 139064
rect 1479 139125 1550 146370
rect 1756 146341 1822 146344
rect 1479 139069 1486 139125
rect 1542 139069 1550 139125
rect 1479 139050 1550 139069
rect 1753 146278 1822 146341
rect -150 135921 -74 135932
rect -150 135865 -140 135921
rect -84 135865 -74 135921
rect -150 135856 -74 135865
rect 1753 135921 1819 146278
rect 1753 135865 1758 135921
rect 1814 135865 1819 135921
rect 1753 135860 1819 135865
rect 1758 135856 1814 135860
rect -144 132659 -60 132668
rect -144 132593 -135 132659
rect -69 132593 -60 132659
rect -144 132582 -60 132593
rect 2020 132649 2086 146250
rect 2020 132584 2086 132593
rect 2284 131159 2350 146156
rect 2279 131099 2350 131159
rect 2554 131145 2621 146069
rect 2819 145902 2893 145958
rect -128 129425 -44 129434
rect -128 129359 -119 129425
rect -53 129359 -44 129425
rect 2279 129420 2345 131099
rect 2279 129364 2284 129420
rect 2340 129364 2345 129420
rect 2279 129359 2345 129364
rect 2533 131049 2621 131145
rect -128 129350 -44 129359
rect 2284 129355 2340 129359
rect -144 126183 -60 126192
rect -144 126117 -139 126183
rect -73 126117 -60 126183
rect -144 126108 -60 126117
rect 2533 126173 2599 131049
rect 2837 130831 2893 145902
rect 2533 126117 2538 126173
rect 2594 126117 2599 126173
rect 2533 126112 2599 126117
rect 2538 126108 2594 126112
rect -166 122951 -82 122960
rect -166 122885 -157 122951
rect -91 122885 -82 122951
rect 2829 122946 2895 130831
rect 2829 122890 2834 122946
rect 2890 122890 2895 122946
rect 2829 122885 2895 122890
rect -166 122876 -82 122885
rect 2834 122881 2890 122885
rect -397 120191 -331 120301
rect -518 120125 -331 120191
rect -518 119540 -452 120125
rect -532 119534 -438 119540
rect -532 119456 -524 119534
rect -446 119456 -438 119534
rect -532 119450 -438 119456
rect -643 118761 -637 118827
rect -571 118761 -289 118827
rect -626 118425 -546 118432
rect -626 118359 -619 118425
rect -553 118359 -546 118425
rect -626 118352 -546 118359
rect -644 118191 -564 118198
rect -644 118125 -637 118191
rect -571 118125 -564 118191
rect -644 118118 -564 118125
rect -634 117811 -538 117818
rect -634 117729 -627 117811
rect -545 117729 -538 117811
rect -634 117722 -538 117729
rect -355 117376 -289 118761
rect -483 117310 -477 117376
rect -411 117310 -289 117376
rect -414 114390 -336 114400
rect -414 114316 -402 114390
rect -346 114316 -336 114390
rect -414 114302 -336 114316
rect -410 111123 -330 111132
rect -410 111057 -401 111123
rect -335 111057 -330 111123
rect -410 111048 -330 111057
rect -406 107894 -332 107904
rect -406 107814 -394 107894
rect -338 107814 -332 107894
rect -406 107802 -332 107814
rect -398 105166 -334 105238
<< via2 >>
rect -465 145561 -409 145627
rect 962 145566 1018 145622
rect -161 142319 -95 142385
rect 1225 142324 1286 142381
rect -172 139069 -116 139125
rect 1486 139069 1542 139125
rect -140 135919 -84 135921
rect -140 135867 -138 135919
rect -138 135867 -86 135919
rect -86 135867 -84 135919
rect -140 135865 -84 135867
rect 1758 135865 1814 135921
rect -135 132593 -69 132659
rect 2020 132593 2086 132649
rect -119 129359 -53 129425
rect 2284 129364 2340 129420
rect -139 126117 -73 126173
rect 2538 126117 2594 126173
rect -157 122885 -91 122951
rect 2834 122890 2890 122946
rect -614 118364 -558 118420
rect -632 118130 -576 118186
rect -622 117734 -550 117806
rect -402 114316 -398 114390
rect -398 114316 -346 114390
rect -401 111057 -335 111123
rect -394 107814 -338 107894
<< metal3 >>
rect -470 145627 -404 145632
rect -470 145561 -465 145627
rect -409 145622 1028 145627
rect -409 145566 962 145622
rect 1018 145566 1028 145622
rect -409 145561 1028 145566
rect -470 145556 -404 145561
rect -166 142385 -90 142390
rect 851 142385 1292 142386
rect -166 142319 -161 142385
rect -95 142381 1292 142385
rect -95 142324 1225 142381
rect 1286 142324 1292 142381
rect -95 142319 1292 142324
rect -166 142314 -90 142319
rect -181 139125 1547 139130
rect -181 139069 -172 139125
rect -116 139069 1486 139125
rect 1542 139069 1547 139125
rect -181 139064 1547 139069
rect -145 135923 -79 135926
rect 1477 135923 1819 135926
rect -145 135921 1819 135923
rect -145 135865 -140 135921
rect -84 135865 1758 135921
rect 1814 135865 1819 135921
rect -145 135863 1819 135865
rect -145 135860 -79 135863
rect 1477 135860 1819 135863
rect -140 132659 -64 132664
rect -140 132593 -135 132659
rect -69 132654 803 132659
rect -69 132649 2091 132654
rect -69 132593 2020 132649
rect 2086 132593 2091 132649
rect -140 132588 -64 132593
rect 621 132588 2091 132593
rect -124 129425 -48 129430
rect -124 129359 -119 129425
rect -53 129420 2345 129425
rect -53 129364 2284 129420
rect 2340 129364 2345 129420
rect -53 129359 2345 129364
rect -124 129354 -48 129359
rect -144 126173 2599 126178
rect -144 126117 -139 126173
rect -73 126117 2538 126173
rect 2594 126117 2599 126173
rect -144 126112 2599 126117
rect -162 122951 -86 122956
rect -162 122885 -157 122951
rect -91 122946 2895 122951
rect -91 122890 2834 122946
rect 2890 122890 2895 122946
rect -91 122885 2895 122890
rect -162 122880 -86 122885
rect -540 118425 -335 118431
rect -619 118420 -335 118425
rect -619 118364 -614 118420
rect -558 118365 -335 118420
rect -558 118364 -540 118365
rect -619 118359 -540 118364
rect -881 118186 -571 118191
rect -881 118130 -632 118186
rect -576 118130 -571 118186
rect -881 118125 -571 118130
rect -881 111123 -815 118125
rect -717 117806 -545 117811
rect -717 117734 -622 117806
rect -550 117734 -545 117806
rect -717 117729 -545 117734
rect -717 111406 -635 117729
rect -401 114400 -335 118365
rect -414 114390 -335 114400
rect -414 114316 -402 114390
rect -346 114374 -335 114390
rect -346 114316 -336 114374
rect -414 114302 -336 114316
rect -722 111326 -716 111406
rect -636 111326 -630 111406
rect -717 111325 -635 111326
rect -406 111123 -330 111128
rect -881 111057 -401 111123
rect -335 111057 -330 111123
rect -406 111052 -330 111057
rect -717 110855 -635 110861
rect -717 107895 -635 110775
rect -406 107900 -332 107904
rect -410 107895 -328 107900
rect -717 107894 -328 107895
rect -717 107814 -394 107894
rect -338 107814 -328 107894
rect -717 107813 -328 107814
rect -410 107802 -328 107813
<< via3 >>
rect -716 111326 -636 111406
rect -717 110775 -635 110855
<< metal4 >>
rect -717 111406 -635 111407
rect -717 111326 -716 111406
rect -636 111326 -635 111406
rect -717 110856 -635 111326
rect -718 110855 -634 110856
rect -718 110775 -717 110855
rect -635 110775 -634 110855
rect -718 110774 -634 110775
use counter_4  counter_4_0
timestamp 1745485683
transform 0 -1 -40 1 0 105408
box -318 0 12226 976
use counter_8  counter_8_0
timestamp 1745486774
transform 0 -1 -40 1 0 120476
box -318 0 25180 976
use decoder_8  decoder_8_0
timestamp 1745492145
transform 1 0 238 0 1 145618
box -238 -145618 5702 1196
use inv  inv_0 ~/magic/library/mag
timestamp 1738780557
transform 0 -1 -40 1 0 119536
box -4 0 322 976
use inv  inv_1
timestamp 1738780557
transform 0 -1 -40 1 0 119844
box -4 0 322 976
use inv  inv_2
timestamp 1738780557
transform 1 0 6572 0 1 -1020
box -4 0 322 976
use inv  inv_3
timestamp 1738780557
transform 1 0 6264 0 1 -1020
box -4 0 322 976
use inv  inv_4
timestamp 1738780557
transform 1 0 7188 0 1 -1020
box -4 0 322 976
use inv  inv_5
timestamp 1738780557
transform 1 0 6880 0 1 -1020
box -4 0 322 976
use inv  inv_6
timestamp 1738780557
transform 1 0 5648 0 1 -1020
box -4 0 322 976
use inv  inv_7
timestamp 1738780557
transform 1 0 5956 0 1 -1020
box -4 0 322 976
use inv  inv_8
timestamp 1738780557
transform 1 0 7804 0 1 -1020
box -4 0 322 976
use inv  inv_9
timestamp 1738780557
transform 1 0 7496 0 1 -1020
box -4 0 322 976
use memory_8  memory_8_0
timestamp 1744679307
transform 1 0 6108 0 1 145480
box -134 -145474 1992 600
use mux4  mux4_0
timestamp 1745483395
transform 0 -1 -40 1 0 117626
box 0 0 1914 976
<< labels >>
flabel metal1 -202 119384 -137 119506 0 FreeSerif 160 270 0 0 Freq1
port 3 nsew
flabel metal2 -398 105166 -334 105238 0 FreeSerif 160 270 0 0 CLK
port 1 nsew
flabel metal1 -963 119428 -898 119550 0 FreeSerif 160 270 0 0 Freq0
port 2 nsew
flabel metal2 436 146748 502 146814 0 FreeSerif 160 0 0 0 Wave1
port 21 nsew
flabel metal2 700 146654 766 146720 0 FreeSerif 160 0 0 0 Wave0
port 20 nsew
flabel locali 5828 -674 5894 -472 0 FreeSerif 160 0 0 0 Y7
port 19 nsew
flabel locali 6136 -674 6202 -472 0 FreeSerif 160 0 0 0 Y6
port 18 nsew
flabel locali 6444 -674 6510 -472 0 FreeSerif 160 0 0 0 Y5
port 17 nsew
flabel locali 6752 -564 6818 -362 0 FreeSerif 160 0 0 0 Y4
port 16 nsew
flabel locali 7060 -584 7126 -382 0 FreeSerif 160 0 0 0 Y3
port 15 nsew
flabel locali 7368 -592 7434 -390 0 FreeSerif 160 0 0 0 Y2
port 14 nsew
flabel locali 7676 -594 7742 -392 0 FreeSerif 160 0 0 0 Y1
port 13 nsew
flabel locali 7984 -598 8050 -396 0 FreeSerif 160 0 0 0 Y0
port 12 nsew
<< end >>
