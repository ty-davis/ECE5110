magic
tech sky130A
timestamp 1744679307
<< nwell >>
rect -27 120 973 300
<< nmos >>
<< pmos >>
<< ndiff >>
rect 581 -1955 614 -1922
rect 614 -1955 706 -1922
rect 332 -1955 365 -1922
rect 116 -1955 208 -1922
rect 863 -1955 955 -1922
rect 489 -1955 581 -1922
rect 738 -1955 830 -1922
rect 365 -1955 457 -1922
rect 240 -1955 332 -1922
rect 83 -1955 116 -1922
rect -9 -1955 83 -1922
rect 830 -1955 863 -1922
rect 581 -2189 614 -2156
rect 614 -2189 706 -2156
rect 332 -2189 365 -2156
rect 116 -2189 208 -2156
rect 863 -2189 955 -2156
rect 489 -2189 581 -2156
rect 738 -2189 830 -2156
rect 365 -2189 457 -2156
rect 240 -2189 332 -2156
rect 83 -2189 116 -2156
rect -9 -2189 83 -2156
rect 830 -2189 863 -2156
rect 581 -2423 614 -2390
rect 614 -2423 706 -2390
rect 332 -2423 365 -2390
rect 116 -2423 208 -2390
rect 863 -2423 955 -2390
rect 489 -2423 581 -2390
rect 738 -2423 830 -2390
rect 365 -2423 457 -2390
rect 240 -2423 332 -2390
rect 83 -2423 116 -2390
rect -9 -2423 83 -2390
rect 830 -2423 863 -2390
rect 581 -2657 614 -2624
rect 614 -2657 706 -2624
rect 332 -2657 365 -2624
rect 116 -2657 208 -2624
rect 863 -2657 955 -2624
rect 489 -2657 581 -2624
rect 738 -2657 830 -2624
rect 365 -2657 457 -2624
rect 240 -2657 332 -2624
rect 83 -2657 116 -2624
rect -9 -2657 83 -2624
rect 830 -2657 863 -2624
rect 581 -2891 614 -2858
rect 614 -2891 706 -2858
rect 332 -2891 365 -2858
rect 116 -2891 208 -2858
rect 863 -2891 955 -2858
rect 489 -2891 581 -2858
rect 738 -2891 830 -2858
rect 365 -2891 457 -2858
rect 240 -2891 332 -2858
rect 83 -2891 116 -2858
rect -9 -2891 83 -2858
rect 830 -2891 863 -2858
rect 581 -3125 614 -3092
rect 614 -3125 706 -3092
rect 332 -3125 365 -3092
rect 116 -3125 208 -3092
rect 863 -3125 955 -3092
rect 489 -3125 581 -3092
rect 738 -3125 830 -3092
rect 365 -3125 457 -3092
rect 240 -3125 332 -3092
rect 83 -3125 116 -3092
rect -9 -3125 83 -3092
rect 830 -3125 863 -3092
rect 581 -3359 614 -3326
rect 614 -3359 706 -3326
rect 332 -3359 365 -3326
rect 116 -3359 208 -3326
rect 863 -3359 955 -3326
rect 489 -3359 581 -3326
rect 738 -3359 830 -3326
rect 365 -3359 457 -3326
rect 240 -3359 332 -3326
rect 83 -3359 116 -3326
rect -9 -3359 83 -3326
rect 830 -3359 863 -3326
rect 581 -3593 614 -3560
rect 614 -3593 706 -3560
rect 332 -3593 365 -3560
rect 116 -3593 208 -3560
rect 863 -3593 955 -3560
rect 489 -3593 581 -3560
rect 738 -3593 830 -3560
rect 365 -3593 457 -3560
rect 240 -3593 332 -3560
rect 83 -3593 116 -3560
rect -9 -3593 83 -3560
rect 830 -3593 863 -3560
rect 581 -3827 614 -3794
rect 614 -3827 706 -3794
rect 863 -3827 955 -3794
rect 489 -3827 581 -3794
rect 738 -3827 830 -3794
rect 830 -3827 863 -3794
rect 581 -4061 614 -4028
rect 614 -4061 706 -4028
rect 332 -4061 365 -4028
rect 863 -4061 955 -4028
rect 489 -4061 581 -4028
rect 738 -4061 830 -4028
rect 365 -4061 457 -4028
rect 240 -4061 332 -4028
rect 830 -4061 863 -4028
rect 581 -4295 614 -4262
rect 614 -4295 706 -4262
rect 332 -4295 365 -4262
rect 116 -4295 208 -4262
rect 863 -4295 955 -4262
rect 489 -4295 581 -4262
rect 738 -4295 830 -4262
rect 365 -4295 457 -4262
rect 240 -4295 332 -4262
rect 83 -4295 116 -4262
rect 830 -4295 863 -4262
rect 581 -4529 614 -4496
rect 614 -4529 706 -4496
rect 332 -4529 365 -4496
rect 116 -4529 208 -4496
rect 863 -4529 955 -4496
rect 489 -4529 581 -4496
rect 738 -4529 830 -4496
rect 365 -4529 457 -4496
rect 83 -4529 116 -4496
rect 240 -4529 332 -4496
rect 830 -4529 863 -4496
rect 581 -4763 614 -4730
rect 614 -4763 706 -4730
rect 332 -4763 365 -4730
rect 116 -4763 208 -4730
rect 863 -4763 955 -4730
rect 489 -4763 581 -4730
rect 738 -4763 830 -4730
rect 365 -4763 457 -4730
rect 240 -4763 332 -4730
rect 83 -4763 116 -4730
rect -9 -4763 83 -4730
rect 830 -4763 863 -4730
rect 581 -4997 614 -4964
rect 614 -4997 706 -4964
rect 332 -4997 365 -4964
rect 863 -4997 955 -4964
rect 489 -4997 581 -4964
rect 738 -4997 830 -4964
rect 365 -4997 457 -4964
rect 83 -4997 116 -4964
rect -9 -4997 83 -4964
rect 240 -4997 332 -4964
rect 830 -4997 863 -4964
rect 581 -5231 614 -5198
rect 614 -5231 706 -5198
rect 332 -5231 365 -5198
rect 116 -5231 208 -5198
rect 863 -5231 955 -5198
rect 489 -5231 581 -5198
rect 738 -5231 830 -5198
rect 365 -5231 457 -5198
rect 240 -5231 332 -5198
rect 83 -5231 116 -5198
rect -9 -5231 83 -5198
rect 830 -5231 863 -5198
rect 581 -5465 614 -5432
rect 614 -5465 706 -5432
rect 332 -5465 365 -5432
rect 116 -5465 208 -5432
rect 863 -5465 955 -5432
rect 489 -5465 581 -5432
rect 738 -5465 830 -5432
rect 365 -5465 457 -5432
rect 83 -5465 116 -5432
rect -9 -5465 83 -5432
rect 240 -5465 332 -5432
rect 830 -5465 863 -5432
rect 581 -5699 614 -5666
rect 614 -5699 706 -5666
rect 332 -5699 365 -5666
rect 116 -5699 208 -5666
rect 863 -5699 955 -5666
rect 489 -5699 581 -5666
rect 738 -5699 830 -5666
rect 365 -5699 457 -5666
rect 240 -5699 332 -5666
rect 83 -5699 116 -5666
rect -9 -5699 83 -5666
rect 830 -5699 863 -5666
rect 581 -5933 614 -5900
rect 614 -5933 706 -5900
rect 332 -5933 365 -5900
rect 116 -5933 208 -5900
rect 863 -5933 955 -5900
rect 489 -5933 581 -5900
rect 738 -5933 830 -5900
rect 365 -5933 457 -5900
rect 83 -5933 116 -5900
rect -9 -5933 83 -5900
rect 830 -5933 863 -5900
rect 581 -6167 614 -6134
rect 614 -6167 706 -6134
rect 332 -6167 365 -6134
rect 863 -6167 955 -6134
rect 489 -6167 581 -6134
rect 738 -6167 830 -6134
rect 365 -6167 457 -6134
rect 240 -6167 332 -6134
rect 83 -6167 116 -6134
rect -9 -6167 83 -6134
rect 830 -6167 863 -6134
rect 581 -6401 614 -6368
rect 614 -6401 706 -6368
rect 332 -6401 365 -6368
rect 863 -6401 955 -6368
rect 489 -6401 581 -6368
rect 738 -6401 830 -6368
rect 365 -6401 457 -6368
rect 83 -6401 116 -6368
rect -9 -6401 83 -6368
rect 830 -6401 863 -6368
rect 581 -6635 614 -6602
rect 614 -6635 706 -6602
rect 332 -6635 365 -6602
rect 116 -6635 208 -6602
rect 863 -6635 955 -6602
rect 489 -6635 581 -6602
rect 738 -6635 830 -6602
rect 365 -6635 457 -6602
rect 240 -6635 332 -6602
rect 83 -6635 116 -6602
rect 830 -6635 863 -6602
rect 581 -6869 614 -6836
rect 614 -6869 706 -6836
rect 332 -6869 365 -6836
rect 116 -6869 208 -6836
rect 863 -6869 955 -6836
rect 489 -6869 581 -6836
rect 738 -6869 830 -6836
rect 365 -6869 457 -6836
rect 83 -6869 116 -6836
rect 830 -6869 863 -6836
rect 581 -7103 614 -7070
rect 614 -7103 706 -7070
rect 332 -7103 365 -7070
rect 863 -7103 955 -7070
rect 489 -7103 581 -7070
rect 738 -7103 830 -7070
rect 365 -7103 457 -7070
rect 240 -7103 332 -7070
rect 830 -7103 863 -7070
rect 581 -7337 614 -7304
rect 614 -7337 706 -7304
rect 332 -7337 365 -7304
rect 863 -7337 955 -7304
rect 489 -7337 581 -7304
rect 738 -7337 830 -7304
rect 365 -7337 457 -7304
rect 830 -7337 863 -7304
rect 581 -7571 614 -7538
rect 614 -7571 706 -7538
rect 863 -7571 955 -7538
rect 738 -7571 830 -7538
rect 830 -7571 863 -7538
rect 581 -7805 614 -7772
rect 614 -7805 706 -7772
rect 332 -7805 365 -7772
rect 863 -7805 955 -7772
rect 489 -7805 581 -7772
rect 738 -7805 830 -7772
rect 365 -7805 457 -7772
rect 830 -7805 863 -7772
rect 581 -8039 614 -8006
rect 614 -8039 706 -8006
rect 332 -8039 365 -8006
rect 863 -8039 955 -8006
rect 489 -8039 581 -8006
rect 738 -8039 830 -8006
rect 365 -8039 457 -8006
rect 240 -8039 332 -8006
rect 830 -8039 863 -8006
rect 581 -8273 614 -8240
rect 614 -8273 706 -8240
rect 332 -8273 365 -8240
rect 863 -8273 955 -8240
rect 489 -8273 581 -8240
rect 738 -8273 830 -8240
rect 240 -8273 332 -8240
rect 365 -8273 457 -8240
rect 830 -8273 863 -8240
rect 581 -8507 614 -8474
rect 614 -8507 706 -8474
rect 332 -8507 365 -8474
rect 116 -8507 208 -8474
rect 863 -8507 955 -8474
rect 489 -8507 581 -8474
rect 738 -8507 830 -8474
rect 365 -8507 457 -8474
rect 240 -8507 332 -8474
rect 83 -8507 116 -8474
rect 830 -8507 863 -8474
rect 581 -8741 614 -8708
rect 614 -8741 706 -8708
rect 332 -8741 365 -8708
rect 116 -8741 208 -8708
rect 863 -8741 955 -8708
rect 489 -8741 581 -8708
rect 738 -8741 830 -8708
rect 83 -8741 116 -8708
rect 365 -8741 457 -8708
rect 830 -8741 863 -8708
rect 581 -8975 614 -8942
rect 614 -8975 706 -8942
rect 332 -8975 365 -8942
rect 116 -8975 208 -8942
rect 863 -8975 955 -8942
rect 489 -8975 581 -8942
rect 738 -8975 830 -8942
rect 365 -8975 457 -8942
rect 83 -8975 116 -8942
rect 240 -8975 332 -8942
rect 830 -8975 863 -8942
rect 581 -9209 614 -9176
rect 614 -9209 706 -9176
rect 332 -9209 365 -9176
rect 116 -9209 208 -9176
rect 863 -9209 955 -9176
rect 489 -9209 581 -9176
rect 738 -9209 830 -9176
rect 240 -9209 332 -9176
rect 83 -9209 116 -9176
rect 365 -9209 457 -9176
rect 830 -9209 863 -9176
rect 581 -9443 614 -9410
rect 614 -9443 706 -9410
rect 332 -9443 365 -9410
rect 116 -9443 208 -9410
rect 863 -9443 955 -9410
rect 489 -9443 581 -9410
rect 738 -9443 830 -9410
rect 365 -9443 457 -9410
rect 240 -9443 332 -9410
rect 83 -9443 116 -9410
rect -9 -9443 83 -9410
rect 830 -9443 863 -9410
rect 581 -9677 614 -9644
rect 614 -9677 706 -9644
rect 332 -9677 365 -9644
rect 863 -9677 955 -9644
rect 489 -9677 581 -9644
rect 738 -9677 830 -9644
rect 83 -9677 116 -9644
rect 365 -9677 457 -9644
rect -9 -9677 83 -9644
rect 830 -9677 863 -9644
rect 581 -9911 614 -9878
rect 614 -9911 706 -9878
rect 332 -9911 365 -9878
rect 863 -9911 955 -9878
rect 489 -9911 581 -9878
rect 738 -9911 830 -9878
rect 365 -9911 457 -9878
rect 83 -9911 116 -9878
rect -9 -9911 83 -9878
rect 240 -9911 332 -9878
rect 830 -9911 863 -9878
rect 581 -10145 614 -10112
rect 614 -10145 706 -10112
rect 332 -10145 365 -10112
rect 863 -10145 955 -10112
rect 489 -10145 581 -10112
rect 738 -10145 830 -10112
rect 240 -10145 332 -10112
rect 83 -10145 116 -10112
rect -9 -10145 83 -10112
rect 365 -10145 457 -10112
rect 830 -10145 863 -10112
rect 581 -10379 614 -10346
rect 614 -10379 706 -10346
rect 332 -10379 365 -10346
rect 116 -10379 208 -10346
rect 863 -10379 955 -10346
rect 489 -10379 581 -10346
rect 738 -10379 830 -10346
rect 365 -10379 457 -10346
rect 240 -10379 332 -10346
rect 83 -10379 116 -10346
rect -9 -10379 83 -10346
rect 830 -10379 863 -10346
rect 581 -10613 614 -10580
rect 614 -10613 706 -10580
rect 332 -10613 365 -10580
rect 116 -10613 208 -10580
rect 863 -10613 955 -10580
rect 489 -10613 581 -10580
rect 738 -10613 830 -10580
rect 83 -10613 116 -10580
rect 365 -10613 457 -10580
rect -9 -10613 83 -10580
rect 830 -10613 863 -10580
rect 581 -10847 614 -10814
rect 614 -10847 706 -10814
rect 332 -10847 365 -10814
rect 116 -10847 208 -10814
rect 863 -10847 955 -10814
rect 489 -10847 581 -10814
rect 738 -10847 830 -10814
rect 365 -10847 457 -10814
rect 83 -10847 116 -10814
rect -9 -10847 83 -10814
rect 240 -10847 332 -10814
rect 830 -10847 863 -10814
rect 581 -11081 614 -11048
rect 614 -11081 706 -11048
rect 332 -11081 365 -11048
rect 116 -11081 208 -11048
rect 863 -11081 955 -11048
rect 489 -11081 581 -11048
rect 738 -11081 830 -11048
rect 240 -11081 332 -11048
rect 83 -11081 116 -11048
rect -9 -11081 83 -11048
rect 365 -11081 457 -11048
rect 830 -11081 863 -11048
rect 830 -11315 863 -11282
rect 738 -11315 830 -11282
rect 581 -11549 614 -11516
rect 614 -11549 706 -11516
rect 332 -11549 365 -11516
rect 863 -11549 955 -11516
rect 489 -11549 581 -11516
rect 738 -11549 830 -11516
rect 365 -11549 457 -11516
rect 830 -11549 863 -11516
rect 581 -11783 614 -11750
rect 614 -11783 706 -11750
rect 332 -11783 365 -11750
rect 863 -11783 955 -11750
rect 489 -11783 581 -11750
rect 365 -11783 457 -11750
rect 240 -11783 332 -11750
rect 830 -11783 863 -11750
rect 581 -12017 614 -11984
rect 614 -12017 706 -11984
rect 332 -12017 365 -11984
rect 116 -12017 208 -11984
rect 863 -12017 955 -11984
rect 489 -12017 581 -11984
rect 738 -12017 830 -11984
rect 83 -12017 116 -11984
rect 240 -12017 332 -11984
rect 830 -12017 863 -11984
rect 581 -12251 614 -12218
rect 332 -12251 365 -12218
rect 489 -12251 581 -12218
rect 83 -12251 116 -12218
rect 365 -12251 457 -12218
rect -9 -12251 83 -12218
rect 581 -12485 614 -12452
rect 614 -12485 706 -12452
rect 332 -12485 365 -12452
rect 116 -12485 208 -12452
rect 83 -12485 116 -12452
rect 365 -12485 457 -12452
rect 240 -12485 332 -12452
rect 738 -12485 830 -12452
rect -9 -12485 83 -12452
rect 830 -12485 863 -12452
rect 581 -12719 614 -12686
rect 332 -12719 365 -12686
rect 116 -12719 208 -12686
rect 489 -12719 581 -12686
rect 83 -12719 116 -12686
rect 738 -12719 830 -12686
rect 365 -12719 457 -12686
rect 240 -12719 332 -12686
rect -9 -12719 83 -12686
rect 830 -12719 863 -12686
rect 581 -12953 614 -12920
rect 614 -12953 706 -12920
rect 332 -12953 365 -12920
rect 116 -12953 208 -12920
rect 863 -12953 955 -12920
rect 83 -12953 116 -12920
rect 365 -12953 457 -12920
rect 240 -12953 332 -12920
rect 489 -12953 581 -12920
rect -9 -12953 83 -12920
rect 830 -12953 863 -12920
rect 581 -13187 614 -13154
rect 614 -13187 706 -13154
rect 332 -13187 365 -13154
rect 116 -13187 208 -13154
rect 863 -13187 955 -13154
rect 489 -13187 581 -13154
rect 738 -13187 830 -13154
rect 365 -13187 457 -13154
rect 240 -13187 332 -13154
rect 83 -13187 116 -13154
rect -9 -13187 83 -13154
rect 830 -13187 863 -13154
rect 581 -13421 614 -13388
rect 614 -13421 706 -13388
rect 332 -13421 365 -13388
rect 116 -13421 208 -13388
rect 863 -13421 955 -13388
rect 83 -13421 116 -13388
rect 365 -13421 457 -13388
rect 240 -13421 332 -13388
rect 738 -13421 830 -13388
rect -9 -13421 83 -13388
rect 489 -13421 581 -13388
rect 830 -13421 863 -13388
rect 581 -13655 614 -13622
rect 614 -13655 706 -13622
rect 332 -13655 365 -13622
rect 116 -13655 208 -13622
rect 489 -13655 581 -13622
rect 83 -13655 116 -13622
rect 738 -13655 830 -13622
rect 365 -13655 457 -13622
rect -9 -13655 83 -13622
rect 830 -13655 863 -13622
rect 581 -13889 614 -13856
rect 332 -13889 365 -13856
rect 83 -13889 116 -13856
rect 489 -13889 581 -13856
rect 365 -13889 457 -13856
rect 240 -13889 332 -13856
rect -9 -13889 83 -13856
rect 581 -14123 614 -14090
rect 614 -14123 706 -14090
rect 332 -14123 365 -14090
rect 116 -14123 208 -14090
rect 863 -14123 955 -14090
rect 83 -14123 116 -14090
rect 738 -14123 830 -14090
rect 240 -14123 332 -14090
rect -9 -14123 83 -14090
rect 830 -14123 863 -14090
rect 581 -14357 614 -14324
rect 614 -14357 706 -14324
rect 332 -14357 365 -14324
rect 116 -14357 208 -14324
rect 863 -14357 955 -14324
rect 489 -14357 581 -14324
rect 738 -14357 830 -14324
rect 83 -14357 116 -14324
rect 365 -14357 457 -14324
rect 240 -14357 332 -14324
rect 830 -14357 863 -14324
rect 581 -14591 614 -14558
rect 614 -14591 706 -14558
rect 332 -14591 365 -14558
rect 863 -14591 955 -14558
rect 365 -14591 457 -14558
rect 240 -14591 332 -14558
rect 830 -14591 863 -14558
rect 830 -14825 863 -14792
rect 489 -14825 581 -14792
rect 581 -14825 614 -14792
rect 738 -14825 830 -14792
rect 157 -1838 208 -1805
rect 655 -1838 706 -1805
rect 489 -1838 540 -1805
rect 738 -1838 789 -1805
rect 904 -1838 955 -1805
rect 240 -1838 291 -1805
rect -9 -1838 42 -1805
rect 406 -1838 457 -1805
rect 157 -2072 208 -2039
rect 655 -2072 706 -2039
rect 489 -2072 540 -2039
rect 738 -2072 789 -2039
rect 904 -2072 955 -2039
rect 240 -2072 291 -2039
rect -9 -2072 42 -2039
rect 406 -2072 457 -2039
rect 157 -2306 208 -2273
rect 655 -2306 706 -2273
rect 489 -2306 540 -2273
rect 738 -2306 789 -2273
rect 904 -2306 955 -2273
rect 240 -2306 291 -2273
rect -9 -2306 42 -2273
rect 406 -2306 457 -2273
rect 157 -2540 208 -2507
rect 655 -2540 706 -2507
rect 489 -2540 540 -2507
rect 738 -2540 789 -2507
rect 904 -2540 955 -2507
rect 240 -2540 291 -2507
rect -9 -2540 42 -2507
rect 406 -2540 457 -2507
rect 157 -2774 208 -2741
rect 655 -2774 706 -2741
rect 489 -2774 540 -2741
rect 738 -2774 789 -2741
rect 904 -2774 955 -2741
rect 240 -2774 291 -2741
rect -9 -2774 42 -2741
rect 406 -2774 457 -2741
rect 157 -3008 208 -2975
rect 655 -3008 706 -2975
rect 489 -3008 540 -2975
rect 738 -3008 789 -2975
rect 904 -3008 955 -2975
rect 240 -3008 291 -2975
rect -9 -3008 42 -2975
rect 406 -3008 457 -2975
rect 157 -3242 208 -3209
rect 655 -3242 706 -3209
rect 489 -3242 540 -3209
rect 738 -3242 789 -3209
rect 904 -3242 955 -3209
rect 240 -3242 291 -3209
rect -9 -3242 42 -3209
rect 406 -3242 457 -3209
rect 157 -3476 208 -3443
rect 655 -3476 706 -3443
rect 489 -3476 540 -3443
rect 738 -3476 789 -3443
rect 904 -3476 955 -3443
rect 240 -3476 291 -3443
rect -9 -3476 42 -3443
rect 406 -3476 457 -3443
rect 157 -3710 208 -3677
rect 655 -3710 706 -3677
rect 489 -3710 540 -3677
rect 738 -3710 789 -3677
rect 904 -3710 955 -3677
rect 240 -3710 291 -3677
rect -9 -3710 42 -3677
rect 406 -3710 457 -3677
rect 655 -3944 706 -3911
rect 489 -3944 540 -3911
rect 738 -3944 789 -3911
rect 904 -3944 955 -3911
rect 406 -3944 457 -3911
rect 655 -4178 706 -4145
rect 489 -4178 540 -4145
rect 738 -4178 789 -4145
rect 904 -4178 955 -4145
rect 240 -4178 291 -4145
rect 406 -4178 457 -4145
rect 157 -4412 208 -4379
rect 655 -4412 706 -4379
rect 489 -4412 540 -4379
rect 738 -4412 789 -4379
rect 904 -4412 955 -4379
rect 406 -4412 457 -4379
rect 157 -4646 208 -4613
rect 655 -4646 706 -4613
rect 489 -4646 540 -4613
rect 738 -4646 789 -4613
rect 904 -4646 955 -4613
rect 240 -4646 291 -4613
rect 406 -4646 457 -4613
rect 655 -4880 706 -4847
rect 489 -4880 540 -4847
rect 738 -4880 789 -4847
rect 904 -4880 955 -4847
rect -9 -4880 42 -4847
rect 406 -4880 457 -4847
rect 655 -5114 706 -5081
rect 489 -5114 540 -5081
rect 738 -5114 789 -5081
rect 904 -5114 955 -5081
rect 240 -5114 291 -5081
rect -9 -5114 42 -5081
rect 406 -5114 457 -5081
rect 157 -5348 208 -5315
rect 655 -5348 706 -5315
rect 489 -5348 540 -5315
rect 738 -5348 789 -5315
rect 904 -5348 955 -5315
rect -9 -5348 42 -5315
rect 406 -5348 457 -5315
rect 157 -5582 208 -5549
rect 655 -5582 706 -5549
rect 489 -5582 540 -5549
rect 738 -5582 789 -5549
rect 904 -5582 955 -5549
rect 240 -5582 291 -5549
rect -9 -5582 42 -5549
rect 406 -5582 457 -5549
rect 157 -5816 208 -5783
rect 655 -5816 706 -5783
rect 489 -5816 540 -5783
rect 738 -5816 789 -5783
rect 904 -5816 955 -5783
rect 240 -5816 291 -5783
rect -9 -5816 42 -5783
rect 406 -5816 457 -5783
rect 157 -6050 208 -6017
rect 655 -6050 706 -6017
rect 489 -6050 540 -6017
rect 738 -6050 789 -6017
rect 904 -6050 955 -6017
rect 240 -6050 291 -6017
rect -9 -6050 42 -6017
rect 406 -6050 457 -6017
rect 655 -6284 706 -6251
rect 489 -6284 540 -6251
rect 738 -6284 789 -6251
rect 904 -6284 955 -6251
rect 240 -6284 291 -6251
rect -9 -6284 42 -6251
rect 406 -6284 457 -6251
rect 157 -6518 208 -6485
rect 655 -6518 706 -6485
rect 489 -6518 540 -6485
rect 738 -6518 789 -6485
rect 904 -6518 955 -6485
rect 240 -6518 291 -6485
rect -9 -6518 42 -6485
rect 406 -6518 457 -6485
rect 157 -6752 208 -6719
rect 655 -6752 706 -6719
rect 489 -6752 540 -6719
rect 738 -6752 789 -6719
rect 904 -6752 955 -6719
rect 240 -6752 291 -6719
rect 406 -6752 457 -6719
rect 157 -6986 208 -6953
rect 655 -6986 706 -6953
rect 489 -6986 540 -6953
rect 738 -6986 789 -6953
rect 904 -6986 955 -6953
rect 240 -6986 291 -6953
rect 406 -6986 457 -6953
rect 655 -7220 706 -7187
rect 489 -7220 540 -7187
rect 738 -7220 789 -7187
rect 904 -7220 955 -7187
rect 240 -7220 291 -7187
rect 406 -7220 457 -7187
rect 655 -7454 706 -7421
rect 489 -7454 540 -7421
rect 738 -7454 789 -7421
rect 904 -7454 955 -7421
rect 655 -7688 706 -7655
rect 489 -7688 540 -7655
rect 738 -7688 789 -7655
rect 904 -7688 955 -7655
rect 655 -7922 706 -7889
rect 489 -7922 540 -7889
rect 738 -7922 789 -7889
rect 904 -7922 955 -7889
rect 406 -7922 457 -7889
rect 655 -8156 706 -8123
rect 489 -8156 540 -8123
rect 738 -8156 789 -8123
rect 904 -8156 955 -8123
rect 240 -8156 291 -8123
rect 655 -8390 706 -8357
rect 489 -8390 540 -8357
rect 738 -8390 789 -8357
rect 904 -8390 955 -8357
rect 240 -8390 291 -8357
rect 406 -8390 457 -8357
rect 157 -8624 208 -8591
rect 655 -8624 706 -8591
rect 738 -8624 789 -8591
rect 489 -8624 540 -8591
rect 904 -8624 955 -8591
rect 157 -8858 208 -8825
rect 655 -8858 706 -8825
rect 738 -8858 789 -8825
rect 489 -8858 540 -8825
rect 904 -8858 955 -8825
rect 406 -8858 457 -8825
rect 157 -9092 208 -9059
rect 655 -9092 706 -9059
rect 738 -9092 789 -9059
rect 489 -9092 540 -9059
rect 904 -9092 955 -9059
rect 240 -9092 291 -9059
rect 157 -9326 208 -9293
rect 655 -9326 706 -9293
rect 738 -9326 789 -9293
rect 489 -9326 540 -9293
rect 904 -9326 955 -9293
rect 240 -9326 291 -9293
rect 406 -9326 457 -9293
rect 655 -9560 706 -9527
rect 489 -9560 540 -9527
rect 738 -9560 789 -9527
rect 904 -9560 955 -9527
rect -9 -9560 42 -9527
rect 655 -9794 706 -9761
rect 489 -9794 540 -9761
rect 738 -9794 789 -9761
rect 904 -9794 955 -9761
rect -9 -9794 42 -9761
rect 406 -9794 457 -9761
rect 655 -10028 706 -9995
rect 489 -10028 540 -9995
rect 738 -10028 789 -9995
rect 904 -10028 955 -9995
rect 240 -10028 291 -9995
rect -9 -10028 42 -9995
rect 655 -10262 706 -10229
rect 489 -10262 540 -10229
rect 738 -10262 789 -10229
rect 904 -10262 955 -10229
rect 240 -10262 291 -10229
rect -9 -10262 42 -10229
rect 406 -10262 457 -10229
rect 157 -10496 208 -10463
rect 655 -10496 706 -10463
rect 738 -10496 789 -10463
rect 489 -10496 540 -10463
rect 904 -10496 955 -10463
rect -9 -10496 42 -10463
rect 157 -10730 208 -10697
rect 655 -10730 706 -10697
rect 738 -10730 789 -10697
rect 489 -10730 540 -10697
rect 904 -10730 955 -10697
rect -9 -10730 42 -10697
rect 406 -10730 457 -10697
rect 157 -10964 208 -10931
rect 655 -10964 706 -10931
rect 738 -10964 789 -10931
rect 489 -10964 540 -10931
rect 904 -10964 955 -10931
rect 240 -10964 291 -10931
rect -9 -10964 42 -10931
rect 157 -11198 208 -11165
rect 655 -11198 706 -11165
rect 738 -11198 789 -11165
rect 904 -11198 955 -11165
rect 240 -11198 291 -11165
rect -9 -11198 42 -11165
rect 406 -11198 457 -11165
rect 489 -11432 540 -11399
rect 738 -11432 789 -11399
rect 655 -11666 706 -11633
rect 904 -11666 955 -11633
rect 240 -11666 291 -11633
rect 406 -11666 457 -11633
rect 157 -11900 208 -11867
rect 655 -11900 706 -11867
rect 489 -11900 540 -11867
rect 738 -11900 789 -11867
rect 904 -11900 955 -11867
rect 240 -11900 291 -11867
rect 406 -11900 457 -11867
rect 157 -12134 208 -12101
rect 655 -12134 706 -12101
rect 738 -12134 789 -12101
rect 904 -12134 955 -12101
rect 240 -12134 291 -12101
rect -9 -12134 42 -12101
rect 489 -12368 540 -12335
rect 240 -12368 291 -12335
rect -9 -12368 42 -12335
rect 406 -12368 457 -12335
rect 157 -12602 208 -12569
rect 655 -12602 706 -12569
rect 738 -12602 789 -12569
rect 489 -12602 540 -12569
rect -9 -12602 42 -12569
rect 406 -12602 457 -12569
rect 157 -12836 208 -12803
rect 655 -12836 706 -12803
rect 489 -12836 540 -12803
rect 738 -12836 789 -12803
rect 904 -12836 955 -12803
rect 240 -12836 291 -12803
rect -9 -12836 42 -12803
rect 406 -12836 457 -12803
rect 157 -13070 208 -13037
rect 655 -13070 706 -13037
rect 489 -13070 540 -13037
rect 904 -13070 955 -13037
rect 738 -13070 789 -13037
rect 240 -13070 291 -13037
rect -9 -13070 42 -13037
rect 406 -13070 457 -13037
rect 157 -13304 208 -13271
rect 655 -13304 706 -13271
rect 489 -13304 540 -13271
rect 904 -13304 955 -13271
rect 240 -13304 291 -13271
rect -9 -13304 42 -13271
rect 406 -13304 457 -13271
rect 157 -13538 208 -13505
rect 489 -13538 540 -13505
rect 738 -13538 789 -13505
rect 240 -13538 291 -13505
rect -9 -13538 42 -13505
rect 406 -13538 457 -13505
rect 157 -13772 208 -13739
rect 655 -13772 706 -13739
rect 738 -13772 789 -13739
rect 240 -13772 291 -13739
rect -9 -13772 42 -13739
rect 406 -13772 457 -13739
rect 489 -14006 540 -13973
rect -9 -14006 42 -13973
rect 406 -14006 457 -13973
rect 157 -14240 208 -14207
rect 655 -14240 706 -14207
rect 738 -14240 789 -14207
rect 489 -14240 540 -14207
rect 904 -14240 955 -14207
rect 240 -14240 291 -14207
rect 655 -14474 706 -14441
rect 489 -14474 540 -14441
rect 904 -14474 955 -14441
rect 240 -14474 291 -14441
rect 406 -14474 457 -14441
rect 655 -14708 706 -14675
rect 489 -14708 540 -14675
rect 738 -14708 789 -14675
rect 904 -14708 955 -14675
rect 406 -14708 457 -14675
rect 738 -14942 789 -14909
rect 904 -10112 955 -10028
rect 904 -2507 955 -2423
rect 904 -2273 955 -2189
rect 904 -12920 955 -12836
rect 904 -4262 955 -4178
rect 904 -6017 955 -5933
rect 904 -3677 955 -3593
rect 904 -10697 955 -10613
rect 904 -7304 955 -7220
rect 904 -3560 955 -3476
rect 904 -8708 955 -8624
rect 904 -10463 955 -10379
rect 904 -5783 955 -5699
rect 904 -13154 955 -13070
rect 904 -5198 955 -5114
rect 904 -8825 955 -8741
rect 904 -8474 955 -8390
rect 904 -14558 955 -14474
rect 904 -2156 955 -2072
rect 904 -5900 955 -5816
rect 904 -3443 955 -3359
rect 904 -4028 955 -3944
rect 904 -6602 955 -6518
rect 904 -5549 955 -5465
rect 904 -11048 955 -10964
rect 904 -10931 955 -10847
rect 904 -9761 955 -9677
rect 904 -5432 955 -5348
rect 904 -14441 955 -14357
rect 904 -8123 955 -8039
rect 904 -9527 955 -9443
rect 904 -4496 955 -4412
rect 904 -10814 955 -10730
rect 904 -2858 955 -2774
rect 904 -10580 955 -10496
rect 904 -8942 955 -8858
rect 904 -5315 955 -5231
rect 904 -6251 955 -6167
rect 904 -4145 955 -4061
rect 904 -14324 955 -14240
rect 904 -11165 955 -11081
rect 904 -10346 955 -10262
rect 904 -9176 955 -9092
rect 904 -8591 955 -8507
rect 904 -7187 955 -7103
rect 904 -8240 955 -8156
rect 904 -8006 955 -7922
rect 904 -1922 955 -1838
rect 904 -4613 955 -4529
rect 904 -14675 955 -14591
rect 904 -11750 955 -11666
rect 904 -5666 955 -5582
rect 904 -10229 955 -10145
rect 904 -7421 955 -7337
rect 904 -13037 955 -12953
rect 904 -6368 955 -6284
rect 904 -2039 955 -1955
rect 904 -13388 955 -13304
rect 904 -4379 955 -4295
rect 904 -11633 955 -11549
rect 904 -9059 955 -8975
rect 904 -7655 955 -7571
rect 904 -2390 955 -2306
rect 904 -6134 955 -6050
rect 904 -9995 955 -9911
rect 904 -9878 955 -9794
rect 904 -2624 955 -2540
rect 904 -11867 955 -11783
rect 904 -3326 955 -3242
rect 904 -9293 955 -9209
rect 904 -5081 955 -4997
rect 904 -13271 955 -13187
rect 904 -8357 955 -8273
rect 904 -4730 955 -4646
rect 904 -12101 955 -12017
rect 904 -2975 955 -2891
rect 904 -3911 955 -3827
rect 904 -7889 955 -7805
rect 904 -2741 955 -2657
rect 904 -11984 955 -11900
rect 904 -4964 955 -4880
rect 904 -4847 955 -4763
rect 904 -3209 955 -3125
rect 904 -7070 955 -6986
rect 904 -6719 955 -6635
rect 904 -9410 955 -9326
rect 904 -9644 955 -9560
rect 904 -3092 955 -3008
rect 904 -6836 955 -6752
rect 904 -6953 955 -6869
rect 904 -7772 955 -7688
rect 904 -6485 955 -6401
rect 904 -14207 955 -14123
rect 738 -10112 789 -10028
rect 738 -2507 789 -2423
rect 738 -12569 789 -12485
rect 738 -2273 789 -2189
rect 738 -4262 789 -4178
rect 738 -6017 789 -5933
rect 738 -3677 789 -3593
rect 738 -10697 789 -10613
rect 738 -7304 789 -7220
rect 738 -14792 789 -14708
rect 738 -3560 789 -3476
rect 738 -8708 789 -8624
rect 738 -10463 789 -10379
rect 738 -5783 789 -5699
rect 738 -11399 789 -11315
rect 738 -13154 789 -13070
rect 738 -5198 789 -5114
rect 738 -8825 789 -8741
rect 738 -8474 789 -8390
rect 738 -11516 789 -11432
rect 738 -12686 789 -12602
rect 738 -2156 789 -2072
rect 738 -5900 789 -5816
rect 738 -3443 789 -3359
rect 738 -4028 789 -3944
rect 738 -6602 789 -6518
rect 738 -5549 789 -5465
rect 738 -11048 789 -10964
rect 738 -10931 789 -10847
rect 738 -9761 789 -9677
rect 738 -5432 789 -5348
rect 738 -8123 789 -8039
rect 738 -9527 789 -9443
rect 738 -4496 789 -4412
rect 738 -10814 789 -10730
rect 738 -2858 789 -2774
rect 738 -10580 789 -10496
rect 738 -8942 789 -8858
rect 738 -5315 789 -5231
rect 738 -6251 789 -6167
rect 738 -4145 789 -4061
rect 738 -14324 789 -14240
rect 738 -11165 789 -11081
rect 738 -10346 789 -10262
rect 738 -9176 789 -9092
rect 738 -8591 789 -8507
rect 738 -7187 789 -7103
rect 738 -8240 789 -8156
rect 738 -8006 789 -7922
rect 738 -1922 789 -1838
rect 738 -4613 789 -4529
rect 738 -5666 789 -5582
rect 738 -10229 789 -10145
rect 738 -7421 789 -7337
rect 738 -6368 789 -6284
rect 738 -13622 789 -13538
rect 738 -2039 789 -1955
rect 738 -4379 789 -4295
rect 738 -9059 789 -8975
rect 738 -12803 789 -12719
rect 738 -7655 789 -7571
rect 738 -2390 789 -2306
rect 738 -6134 789 -6050
rect 738 -9995 789 -9911
rect 738 -9878 789 -9794
rect 738 -2624 789 -2540
rect 738 -13505 789 -13421
rect 738 -3326 789 -3242
rect 738 -9293 789 -9209
rect 738 -5081 789 -4997
rect 738 -13739 789 -13655
rect 738 -8357 789 -8273
rect 738 -4730 789 -4646
rect 738 -12101 789 -12017
rect 738 -2975 789 -2891
rect 738 -3911 789 -3827
rect 738 -7889 789 -7805
rect 738 -2741 789 -2657
rect 738 -11984 789 -11900
rect 738 -4964 789 -4880
rect 738 -4847 789 -4763
rect 738 -3209 789 -3125
rect 738 -7070 789 -6986
rect 738 -6719 789 -6635
rect 738 -9410 789 -9326
rect 738 -9644 789 -9560
rect 738 -3092 789 -3008
rect 738 -6836 789 -6752
rect 738 -6953 789 -6869
rect 738 -14909 789 -14825
rect 738 -7772 789 -7688
rect 738 -6485 789 -6401
rect 738 -14207 789 -14123
rect 655 -10112 706 -10028
rect 655 -2507 706 -2423
rect 655 -12569 706 -12485
rect 655 -2273 706 -2189
rect 655 -12920 706 -12836
rect 655 -4262 706 -4178
rect 655 -6017 706 -5933
rect 655 -3677 706 -3593
rect 655 -10697 706 -10613
rect 655 -7304 706 -7220
rect 655 -3560 706 -3476
rect 655 -8708 706 -8624
rect 655 -10463 706 -10379
rect 655 -5783 706 -5699
rect 655 -13154 706 -13070
rect 655 -5198 706 -5114
rect 655 -8825 706 -8741
rect 655 -8474 706 -8390
rect 655 -14558 706 -14474
rect 655 -2156 706 -2072
rect 655 -5900 706 -5816
rect 655 -3443 706 -3359
rect 655 -4028 706 -3944
rect 655 -6602 706 -6518
rect 655 -5549 706 -5465
rect 655 -11048 706 -10964
rect 655 -10931 706 -10847
rect 655 -9761 706 -9677
rect 655 -5432 706 -5348
rect 655 -8123 706 -8039
rect 655 -9527 706 -9443
rect 655 -4496 706 -4412
rect 655 -10814 706 -10730
rect 655 -2858 706 -2774
rect 655 -10580 706 -10496
rect 655 -8942 706 -8858
rect 655 -5315 706 -5231
rect 655 -6251 706 -6167
rect 655 -4145 706 -4061
rect 655 -14324 706 -14240
rect 655 -11165 706 -11081
rect 655 -10346 706 -10262
rect 655 -9176 706 -9092
rect 655 -8591 706 -8507
rect 655 -7187 706 -7103
rect 655 -8240 706 -8156
rect 655 -8006 706 -7922
rect 655 -1922 706 -1838
rect 655 -4613 706 -4529
rect 655 -14675 706 -14591
rect 655 -11750 706 -11666
rect 655 -5666 706 -5582
rect 655 -10229 706 -10145
rect 655 -7421 706 -7337
rect 655 -13037 706 -12953
rect 655 -6368 706 -6284
rect 655 -2039 706 -1955
rect 655 -13388 706 -13304
rect 655 -4379 706 -4295
rect 655 -11633 706 -11549
rect 655 -9059 706 -8975
rect 655 -7655 706 -7571
rect 655 -2390 706 -2306
rect 655 -6134 706 -6050
rect 655 -9995 706 -9911
rect 655 -9878 706 -9794
rect 655 -2624 706 -2540
rect 655 -3326 706 -3242
rect 655 -9293 706 -9209
rect 655 -5081 706 -4997
rect 655 -13271 706 -13187
rect 655 -13739 706 -13655
rect 655 -8357 706 -8273
rect 655 -4730 706 -4646
rect 655 -12101 706 -12017
rect 655 -2975 706 -2891
rect 655 -3911 706 -3827
rect 655 -7889 706 -7805
rect 655 -2741 706 -2657
rect 655 -11984 706 -11900
rect 655 -4964 706 -4880
rect 655 -4847 706 -4763
rect 655 -3209 706 -3125
rect 655 -7070 706 -6986
rect 655 -6719 706 -6635
rect 655 -9410 706 -9326
rect 655 -9644 706 -9560
rect 655 -3092 706 -3008
rect 655 -6836 706 -6752
rect 655 -6953 706 -6869
rect 655 -7772 706 -7688
rect 655 -6485 706 -6401
rect 655 -14207 706 -14123
rect 489 -10112 540 -10028
rect 489 -2507 540 -2423
rect 489 -2273 540 -2189
rect 489 -4262 540 -4178
rect 489 -6017 540 -5933
rect 489 -3677 540 -3593
rect 489 -7304 540 -7220
rect 489 -14792 540 -14708
rect 489 -3560 540 -3476
rect 489 -8708 540 -8624
rect 489 -5783 540 -5699
rect 489 -13154 540 -13070
rect 489 -5198 540 -5114
rect 489 -8474 540 -8390
rect 489 -11516 540 -11432
rect 489 -12686 540 -12602
rect 489 -2156 540 -2072
rect 489 -5900 540 -5816
rect 489 -3443 540 -3359
rect 489 -4028 540 -3944
rect 489 -6602 540 -6518
rect 489 -5549 540 -5465
rect 489 -11048 540 -10964
rect 489 -5432 540 -5348
rect 489 -14441 540 -14357
rect 489 -4496 540 -4412
rect 489 -10814 540 -10730
rect 489 -13973 540 -13889
rect 489 -2858 540 -2774
rect 489 -10580 540 -10496
rect 489 -8942 540 -8858
rect 489 -5315 540 -5231
rect 489 -6251 540 -6167
rect 489 -4145 540 -4061
rect 489 -14324 540 -14240
rect 489 -10346 540 -10262
rect 489 -9176 540 -9092
rect 489 -7187 540 -7103
rect 489 -8240 540 -8156
rect 489 -8006 540 -7922
rect 489 -1922 540 -1838
rect 489 -4613 540 -4529
rect 489 -5666 540 -5582
rect 489 -7421 540 -7337
rect 489 -13037 540 -12953
rect 489 -6368 540 -6284
rect 489 -13622 540 -13538
rect 489 -2039 540 -1955
rect 489 -4379 540 -4295
rect 489 -12803 540 -12719
rect 489 -2390 540 -2306
rect 489 -6134 540 -6050
rect 489 -9878 540 -9794
rect 489 -2624 540 -2540
rect 489 -13505 540 -13421
rect 489 -11867 540 -11783
rect 489 -3326 540 -3242
rect 489 -5081 540 -4997
rect 489 -13271 540 -13187
rect 489 -4730 540 -4646
rect 489 -2975 540 -2891
rect 489 -3911 540 -3827
rect 489 -2741 540 -2657
rect 489 -11984 540 -11900
rect 489 -12335 540 -12251
rect 489 -4964 540 -4880
rect 489 -4847 540 -4763
rect 489 -3209 540 -3125
rect 489 -7070 540 -6986
rect 489 -6719 540 -6635
rect 489 -9410 540 -9326
rect 489 -9644 540 -9560
rect 489 -3092 540 -3008
rect 489 -6836 540 -6752
rect 489 -6953 540 -6869
rect 489 -7772 540 -7688
rect 489 -6485 540 -6401
rect 406 -3326 457 -3242
rect 406 -2507 457 -2423
rect 406 -9293 457 -9209
rect 406 -2156 457 -2072
rect 406 -13271 457 -13187
rect 406 -2273 457 -2189
rect 406 -5900 457 -5816
rect 406 -12920 457 -12836
rect 406 -8006 457 -7922
rect 406 -8357 457 -8273
rect 406 -1922 457 -1838
rect 406 -4730 457 -4646
rect 406 -2975 457 -2891
rect 406 -14675 457 -14591
rect 406 -3443 457 -3359
rect 406 -4262 457 -4178
rect 406 -7889 457 -7805
rect 406 -5666 457 -5582
rect 406 -10229 457 -10145
rect 406 -3677 457 -3593
rect 406 -13037 457 -12953
rect 406 -2741 457 -2657
rect 406 -4028 457 -3944
rect 406 -12335 457 -12251
rect 406 -4964 457 -4880
rect 406 -6368 457 -6284
rect 406 -13622 457 -13538
rect 406 -6602 457 -6518
rect 406 -2039 457 -1955
rect 406 -13388 457 -13304
rect 406 -3209 457 -3125
rect 406 -10697 457 -10613
rect 406 -7304 457 -7220
rect 406 -3560 457 -3476
rect 406 -7070 457 -6986
rect 406 -9761 457 -9677
rect 406 -5432 457 -5348
rect 406 -12452 457 -12368
rect 406 -9410 457 -9326
rect 406 -14441 457 -14357
rect 406 -11633 457 -11549
rect 406 -3092 457 -3008
rect 406 -4496 457 -4412
rect 406 -5198 457 -5114
rect 406 -6836 457 -6752
rect 406 -13154 457 -13070
rect 406 -10814 457 -10730
rect 406 -13973 457 -13889
rect 406 -2858 457 -2774
rect 406 -2390 457 -2306
rect 406 -8825 457 -8741
rect 406 -8942 457 -8858
rect 406 -6134 457 -6050
rect 406 -8474 457 -8390
rect 406 -9878 457 -9794
rect 406 -13856 457 -13772
rect 406 -11165 457 -11081
rect 406 -12686 457 -12602
rect 406 -10346 457 -10262
rect 406 -2624 457 -2540
rect 406 -11867 457 -11783
rect 240 -3326 291 -3242
rect 240 -2507 291 -2423
rect 240 -5081 291 -4997
rect 240 -2156 291 -2072
rect 240 -8240 291 -8156
rect 240 -9293 291 -9209
rect 240 -10112 291 -10028
rect 240 -13271 291 -13187
rect 240 -2273 291 -2189
rect 240 -12920 291 -12836
rect 240 -8357 291 -8273
rect 240 -1922 291 -1838
rect 240 -4613 291 -4529
rect 240 -4730 291 -4646
rect 240 -2975 291 -2891
rect 240 -11867 291 -11783
rect 240 -12101 291 -12017
rect 240 -3443 291 -3359
rect 240 -4262 291 -4178
rect 240 -11750 291 -11666
rect 240 -5666 291 -5582
rect 240 -10229 291 -10145
rect 240 -3677 291 -3593
rect 240 -13037 291 -12953
rect 240 -2741 291 -2657
rect 240 -6602 291 -6518
rect 240 -2039 291 -1955
rect 240 -5549 291 -5465
rect 240 -13388 291 -13304
rect 240 -3209 291 -3125
rect 240 -3560 291 -3476
rect 240 -11048 291 -10964
rect 240 -7070 291 -6986
rect 240 -10931 291 -10847
rect 240 -12452 291 -12368
rect 240 -5783 291 -5699
rect 240 -6719 291 -6635
rect 240 -9410 291 -9326
rect 240 -14441 291 -14357
rect 240 -8123 291 -8039
rect 240 -9059 291 -8975
rect 240 -12803 291 -12719
rect 240 -3092 291 -3008
rect 240 -13154 291 -13070
rect 240 -5198 291 -5114
rect 240 -2858 291 -2774
rect 240 -2390 291 -2306
rect 240 -6134 291 -6050
rect 240 -8474 291 -8390
rect 240 -9995 291 -9911
rect 240 -6251 291 -6167
rect 240 -4145 291 -4061
rect 240 -13856 291 -13772
rect 240 -14558 291 -14474
rect 240 -11165 291 -11081
rect 240 -10346 291 -10262
rect 240 -9176 291 -9092
rect 240 -2624 291 -2540
rect 240 -13505 291 -13421
rect 240 -7187 291 -7103
rect 240 -14207 291 -14123
rect 157 -3326 208 -3242
rect 157 -2507 208 -2423
rect 157 -9293 208 -9209
rect 157 -2156 208 -2072
rect 157 -12569 208 -12485
rect 157 -13271 208 -13187
rect 157 -2273 208 -2189
rect 157 -5900 208 -5816
rect 157 -12920 208 -12836
rect 157 -13739 208 -13655
rect 157 -1922 208 -1838
rect 157 -4613 208 -4529
rect 157 -4730 208 -4646
rect 157 -2975 208 -2891
rect 157 -12101 208 -12017
rect 157 -3443 208 -3359
rect 157 -5666 208 -5582
rect 157 -6017 208 -5933
rect 157 -3677 208 -3593
rect 157 -13037 208 -12953
rect 157 -2741 208 -2657
rect 157 -11984 208 -11900
rect 157 -13622 208 -13538
rect 157 -6602 208 -6518
rect 157 -2039 208 -1955
rect 157 -5549 208 -5465
rect 157 -13388 208 -13304
rect 157 -3209 208 -3125
rect 157 -10697 208 -10613
rect 157 -3560 208 -3476
rect 157 -8708 208 -8624
rect 157 -11048 208 -10964
rect 157 -10931 208 -10847
rect 157 -4379 208 -4295
rect 157 -10463 208 -10379
rect 157 -5432 208 -5348
rect 157 -5783 208 -5699
rect 157 -6719 208 -6635
rect 157 -9410 208 -9326
rect 157 -9059 208 -8975
rect 157 -12803 208 -12719
rect 157 -3092 208 -3008
rect 157 -4496 208 -4412
rect 157 -6836 208 -6752
rect 157 -13154 208 -13070
rect 157 -6953 208 -6869
rect 157 -10814 208 -10730
rect 157 -2858 208 -2774
rect 157 -2390 208 -2306
rect 157 -8825 208 -8741
rect 157 -8942 208 -8858
rect 157 -10580 208 -10496
rect 157 -5315 208 -5231
rect 157 -14324 208 -14240
rect 157 -11165 208 -11081
rect 157 -12686 208 -12602
rect 157 -9176 208 -9092
rect 157 -2624 208 -2540
rect 157 -8591 208 -8507
rect 157 -13505 208 -13421
rect 157 -14207 208 -14123
rect -9 -3326 42 -3242
rect -9 -2507 42 -2423
rect -9 -5081 42 -4997
rect -9 -2156 42 -2072
rect -9 -10112 42 -10028
rect -9 -12569 42 -12485
rect -9 -13271 42 -13187
rect -9 -2273 42 -2189
rect -9 -5900 42 -5816
rect -9 -12920 42 -12836
rect -9 -13739 42 -13655
rect -9 -1922 42 -1838
rect -9 -2975 42 -2891
rect -9 -3443 42 -3359
rect -9 -14090 42 -14006
rect -9 -5666 42 -5582
rect -9 -6017 42 -5933
rect -9 -10229 42 -10145
rect -9 -3677 42 -3593
rect -9 -13037 42 -12953
rect -9 -2741 42 -2657
rect -9 -12218 42 -12134
rect -9 -12335 42 -12251
rect -9 -4964 42 -4880
rect -9 -6368 42 -6284
rect -9 -13622 42 -13538
rect -9 -2039 42 -1955
rect -9 -4847 42 -4763
rect -9 -5549 42 -5465
rect -9 -3209 42 -3125
rect -9 -13388 42 -13304
rect -9 -10697 42 -10613
rect -9 -3560 42 -3476
rect -9 -11048 42 -10964
rect -9 -10931 42 -10847
rect -9 -9761 42 -9677
rect -9 -10463 42 -10379
rect -9 -5432 42 -5348
rect -9 -5783 42 -5699
rect -9 -12452 42 -12368
rect -9 -9527 42 -9443
rect -9 -9644 42 -9560
rect -9 -12803 42 -12719
rect -9 -3092 42 -3008
rect -9 -13154 42 -13070
rect -9 -5198 42 -5114
rect -9 -10814 42 -10730
rect -9 -13973 42 -13889
rect -9 -2858 42 -2774
rect -9 -2390 42 -2306
rect -9 -10580 42 -10496
rect -9 -6134 42 -6050
rect -9 -5315 42 -5231
rect -9 -9995 42 -9911
rect -9 -6251 42 -6167
rect -9 -9878 42 -9794
rect -9 -13856 42 -13772
rect -9 -11165 42 -11081
rect -9 -12686 42 -12602
rect -9 -10346 42 -10262
rect -9 -2624 42 -2540
rect -9 -13505 42 -13421
rect -9 -6485 42 -6401
<< pdiff >>
rect 904 138 955 227
rect 738 138 789 227
rect 655 138 706 227
rect 489 138 540 227
rect 406 138 457 227
rect 240 138 291 227
rect 157 138 208 227
rect -9 138 42 227
<< ndiffc >>
<< pdiffc >>
rect 921 146 938 163
rect 912 202 947 219
rect 755 146 772 163
rect 746 202 781 219
rect 672 146 689 163
rect 663 202 698 219
rect 506 146 523 163
rect 497 202 532 219
rect 423 146 440 163
rect 414 202 449 219
rect 257 146 274 163
rect 248 202 283 219
rect 174 146 191 163
rect 165 202 200 219
rect 8 146 25 163
rect -1 202 34 219
<< psubdiff >>
rect -27 79 973 107
<< nsubdiff >>
rect -9 254 955 282
<< psubdiffcont >>
rect -15 79 961 107
<< nsubdiffcont >>
rect 3 254 943 282
<< ndcontact >>
rect 589 -1947 606 -1930
rect 340 -1947 357 -1930
rect 91 -1947 108 -1930
rect 838 -1947 855 -1930
rect 589 -2181 606 -2164
rect 340 -2181 357 -2164
rect 91 -2181 108 -2164
rect 838 -2181 855 -2164
rect 589 -2415 606 -2398
rect 340 -2415 357 -2398
rect 91 -2415 108 -2398
rect 838 -2415 855 -2398
rect 589 -2649 606 -2632
rect 340 -2649 357 -2632
rect 91 -2649 108 -2632
rect 838 -2649 855 -2632
rect 589 -2883 606 -2866
rect 340 -2883 357 -2866
rect 91 -2883 108 -2866
rect 838 -2883 855 -2866
rect 589 -3117 606 -3100
rect 340 -3117 357 -3100
rect 91 -3117 108 -3100
rect 838 -3117 855 -3100
rect 589 -3351 606 -3334
rect 340 -3351 357 -3334
rect 91 -3351 108 -3334
rect 838 -3351 855 -3334
rect 589 -3585 606 -3568
rect 340 -3585 357 -3568
rect 91 -3585 108 -3568
rect 838 -3585 855 -3568
rect 589 -3819 606 -3802
rect 838 -3819 855 -3802
rect 589 -4053 606 -4036
rect 340 -4053 357 -4036
rect 838 -4053 855 -4036
rect 589 -4287 606 -4270
rect 340 -4287 357 -4270
rect 91 -4287 108 -4270
rect 838 -4287 855 -4270
rect 589 -4521 606 -4504
rect 340 -4521 357 -4504
rect 91 -4521 108 -4504
rect 838 -4521 855 -4504
rect 589 -4755 606 -4738
rect 340 -4755 357 -4738
rect 91 -4755 108 -4738
rect 838 -4755 855 -4738
rect 589 -4989 606 -4972
rect 340 -4989 357 -4972
rect 91 -4989 108 -4972
rect 838 -4989 855 -4972
rect 589 -5223 606 -5206
rect 340 -5223 357 -5206
rect 91 -5223 108 -5206
rect 838 -5223 855 -5206
rect 589 -5457 606 -5440
rect 340 -5457 357 -5440
rect 91 -5457 108 -5440
rect 838 -5457 855 -5440
rect 589 -5691 606 -5674
rect 340 -5691 357 -5674
rect 91 -5691 108 -5674
rect 838 -5691 855 -5674
rect 589 -5925 606 -5908
rect 340 -5925 357 -5908
rect 91 -5925 108 -5908
rect 838 -5925 855 -5908
rect 589 -6159 606 -6142
rect 340 -6159 357 -6142
rect 91 -6159 108 -6142
rect 838 -6159 855 -6142
rect 589 -6393 606 -6376
rect 340 -6393 357 -6376
rect 91 -6393 108 -6376
rect 838 -6393 855 -6376
rect 589 -6627 606 -6610
rect 340 -6627 357 -6610
rect 91 -6627 108 -6610
rect 838 -6627 855 -6610
rect 589 -6861 606 -6844
rect 340 -6861 357 -6844
rect 91 -6861 108 -6844
rect 838 -6861 855 -6844
rect 589 -7095 606 -7078
rect 340 -7095 357 -7078
rect 838 -7095 855 -7078
rect 589 -7329 606 -7312
rect 340 -7329 357 -7312
rect 838 -7329 855 -7312
rect 589 -7563 606 -7546
rect 838 -7563 855 -7546
rect 589 -7797 606 -7780
rect 340 -7797 357 -7780
rect 838 -7797 855 -7780
rect 589 -8031 606 -8014
rect 340 -8031 357 -8014
rect 838 -8031 855 -8014
rect 589 -8265 606 -8248
rect 340 -8265 357 -8248
rect 838 -8265 855 -8248
rect 589 -8499 606 -8482
rect 340 -8499 357 -8482
rect 91 -8499 108 -8482
rect 838 -8499 855 -8482
rect 589 -8733 606 -8716
rect 340 -8733 357 -8716
rect 91 -8733 108 -8716
rect 838 -8733 855 -8716
rect 589 -8967 606 -8950
rect 340 -8967 357 -8950
rect 91 -8967 108 -8950
rect 838 -8967 855 -8950
rect 589 -9201 606 -9184
rect 340 -9201 357 -9184
rect 91 -9201 108 -9184
rect 838 -9201 855 -9184
rect 589 -9435 606 -9418
rect 340 -9435 357 -9418
rect 91 -9435 108 -9418
rect 838 -9435 855 -9418
rect 589 -9669 606 -9652
rect 340 -9669 357 -9652
rect 91 -9669 108 -9652
rect 838 -9669 855 -9652
rect 589 -9903 606 -9886
rect 340 -9903 357 -9886
rect 91 -9903 108 -9886
rect 838 -9903 855 -9886
rect 589 -10137 606 -10120
rect 340 -10137 357 -10120
rect 91 -10137 108 -10120
rect 838 -10137 855 -10120
rect 589 -10371 606 -10354
rect 340 -10371 357 -10354
rect 91 -10371 108 -10354
rect 838 -10371 855 -10354
rect 589 -10605 606 -10588
rect 340 -10605 357 -10588
rect 91 -10605 108 -10588
rect 838 -10605 855 -10588
rect 589 -10839 606 -10822
rect 340 -10839 357 -10822
rect 91 -10839 108 -10822
rect 838 -10839 855 -10822
rect 589 -11073 606 -11056
rect 340 -11073 357 -11056
rect 91 -11073 108 -11056
rect 838 -11073 855 -11056
rect 838 -11307 855 -11290
rect 589 -11541 606 -11524
rect 340 -11541 357 -11524
rect 838 -11541 855 -11524
rect 589 -11775 606 -11758
rect 340 -11775 357 -11758
rect 838 -11775 855 -11758
rect 589 -12009 606 -11992
rect 340 -12009 357 -11992
rect 91 -12009 108 -11992
rect 838 -12009 855 -11992
rect 589 -12243 606 -12226
rect 340 -12243 357 -12226
rect 91 -12243 108 -12226
rect 589 -12477 606 -12460
rect 340 -12477 357 -12460
rect 91 -12477 108 -12460
rect 838 -12477 855 -12460
rect 589 -12711 606 -12694
rect 340 -12711 357 -12694
rect 91 -12711 108 -12694
rect 838 -12711 855 -12694
rect 589 -12945 606 -12928
rect 340 -12945 357 -12928
rect 91 -12945 108 -12928
rect 838 -12945 855 -12928
rect 589 -13179 606 -13162
rect 340 -13179 357 -13162
rect 91 -13179 108 -13162
rect 838 -13179 855 -13162
rect 589 -13413 606 -13396
rect 340 -13413 357 -13396
rect 91 -13413 108 -13396
rect 838 -13413 855 -13396
rect 589 -13647 606 -13630
rect 340 -13647 357 -13630
rect 91 -13647 108 -13630
rect 838 -13647 855 -13630
rect 589 -13881 606 -13864
rect 340 -13881 357 -13864
rect 91 -13881 108 -13864
rect 589 -14115 606 -14098
rect 340 -14115 357 -14098
rect 91 -14115 108 -14098
rect 838 -14115 855 -14098
rect 589 -14349 606 -14332
rect 340 -14349 357 -14332
rect 91 -14349 108 -14332
rect 838 -14349 855 -14332
rect 589 -14583 606 -14566
rect 340 -14583 357 -14566
rect 838 -14583 855 -14566
rect 838 -14817 855 -14800
rect 589 -14817 606 -14800
rect 174 -1830 191 -1813
rect 672 -1830 689 -1813
rect 506 -1830 523 -1813
rect 755 -1830 772 -1813
rect 921 -1830 938 -1813
rect 257 -1830 274 -1813
rect 8 -1830 25 -1813
rect 423 -1830 440 -1813
rect 174 -2064 191 -2047
rect 672 -2064 689 -2047
rect 506 -2064 523 -2047
rect 755 -2064 772 -2047
rect 921 -2064 938 -2047
rect 257 -2064 274 -2047
rect 8 -2064 25 -2047
rect 423 -2064 440 -2047
rect 174 -2298 191 -2281
rect 672 -2298 689 -2281
rect 506 -2298 523 -2281
rect 755 -2298 772 -2281
rect 921 -2298 938 -2281
rect 257 -2298 274 -2281
rect 8 -2298 25 -2281
rect 423 -2298 440 -2281
rect 174 -2532 191 -2515
rect 672 -2532 689 -2515
rect 506 -2532 523 -2515
rect 755 -2532 772 -2515
rect 921 -2532 938 -2515
rect 257 -2532 274 -2515
rect 8 -2532 25 -2515
rect 423 -2532 440 -2515
rect 174 -2766 191 -2749
rect 672 -2766 689 -2749
rect 506 -2766 523 -2749
rect 755 -2766 772 -2749
rect 921 -2766 938 -2749
rect 257 -2766 274 -2749
rect 8 -2766 25 -2749
rect 423 -2766 440 -2749
rect 174 -3000 191 -2983
rect 672 -3000 689 -2983
rect 506 -3000 523 -2983
rect 755 -3000 772 -2983
rect 921 -3000 938 -2983
rect 257 -3000 274 -2983
rect 8 -3000 25 -2983
rect 423 -3000 440 -2983
rect 174 -3234 191 -3217
rect 672 -3234 689 -3217
rect 506 -3234 523 -3217
rect 755 -3234 772 -3217
rect 921 -3234 938 -3217
rect 257 -3234 274 -3217
rect 8 -3234 25 -3217
rect 423 -3234 440 -3217
rect 174 -3468 191 -3451
rect 672 -3468 689 -3451
rect 506 -3468 523 -3451
rect 755 -3468 772 -3451
rect 921 -3468 938 -3451
rect 257 -3468 274 -3451
rect 8 -3468 25 -3451
rect 423 -3468 440 -3451
rect 174 -3702 191 -3685
rect 672 -3702 689 -3685
rect 506 -3702 523 -3685
rect 755 -3702 772 -3685
rect 921 -3702 938 -3685
rect 257 -3702 274 -3685
rect 8 -3702 25 -3685
rect 423 -3702 440 -3685
rect 672 -3936 689 -3919
rect 506 -3936 523 -3919
rect 755 -3936 772 -3919
rect 921 -3936 938 -3919
rect 423 -3936 440 -3919
rect 672 -4170 689 -4153
rect 506 -4170 523 -4153
rect 755 -4170 772 -4153
rect 921 -4170 938 -4153
rect 257 -4170 274 -4153
rect 423 -4170 440 -4153
rect 174 -4404 191 -4387
rect 672 -4404 689 -4387
rect 506 -4404 523 -4387
rect 755 -4404 772 -4387
rect 921 -4404 938 -4387
rect 423 -4404 440 -4387
rect 174 -4638 191 -4621
rect 672 -4638 689 -4621
rect 506 -4638 523 -4621
rect 755 -4638 772 -4621
rect 921 -4638 938 -4621
rect 257 -4638 274 -4621
rect 423 -4638 440 -4621
rect 672 -4872 689 -4855
rect 506 -4872 523 -4855
rect 755 -4872 772 -4855
rect 921 -4872 938 -4855
rect 8 -4872 25 -4855
rect 423 -4872 440 -4855
rect 672 -5106 689 -5089
rect 506 -5106 523 -5089
rect 755 -5106 772 -5089
rect 921 -5106 938 -5089
rect 257 -5106 274 -5089
rect 8 -5106 25 -5089
rect 423 -5106 440 -5089
rect 174 -5340 191 -5323
rect 672 -5340 689 -5323
rect 506 -5340 523 -5323
rect 755 -5340 772 -5323
rect 921 -5340 938 -5323
rect 8 -5340 25 -5323
rect 423 -5340 440 -5323
rect 174 -5574 191 -5557
rect 672 -5574 689 -5557
rect 506 -5574 523 -5557
rect 755 -5574 772 -5557
rect 921 -5574 938 -5557
rect 257 -5574 274 -5557
rect 8 -5574 25 -5557
rect 423 -5574 440 -5557
rect 174 -5808 191 -5791
rect 672 -5808 689 -5791
rect 506 -5808 523 -5791
rect 755 -5808 772 -5791
rect 921 -5808 938 -5791
rect 257 -5808 274 -5791
rect 8 -5808 25 -5791
rect 423 -5808 440 -5791
rect 174 -6042 191 -6025
rect 672 -6042 689 -6025
rect 506 -6042 523 -6025
rect 755 -6042 772 -6025
rect 921 -6042 938 -6025
rect 257 -6042 274 -6025
rect 8 -6042 25 -6025
rect 423 -6042 440 -6025
rect 672 -6276 689 -6259
rect 506 -6276 523 -6259
rect 755 -6276 772 -6259
rect 921 -6276 938 -6259
rect 257 -6276 274 -6259
rect 8 -6276 25 -6259
rect 423 -6276 440 -6259
rect 174 -6510 191 -6493
rect 672 -6510 689 -6493
rect 506 -6510 523 -6493
rect 755 -6510 772 -6493
rect 921 -6510 938 -6493
rect 257 -6510 274 -6493
rect 8 -6510 25 -6493
rect 423 -6510 440 -6493
rect 174 -6744 191 -6727
rect 672 -6744 689 -6727
rect 506 -6744 523 -6727
rect 755 -6744 772 -6727
rect 921 -6744 938 -6727
rect 257 -6744 274 -6727
rect 423 -6744 440 -6727
rect 174 -6978 191 -6961
rect 672 -6978 689 -6961
rect 506 -6978 523 -6961
rect 755 -6978 772 -6961
rect 921 -6978 938 -6961
rect 257 -6978 274 -6961
rect 423 -6978 440 -6961
rect 672 -7212 689 -7195
rect 506 -7212 523 -7195
rect 755 -7212 772 -7195
rect 921 -7212 938 -7195
rect 257 -7212 274 -7195
rect 423 -7212 440 -7195
rect 672 -7446 689 -7429
rect 506 -7446 523 -7429
rect 755 -7446 772 -7429
rect 921 -7446 938 -7429
rect 672 -7680 689 -7663
rect 506 -7680 523 -7663
rect 755 -7680 772 -7663
rect 921 -7680 938 -7663
rect 672 -7914 689 -7897
rect 506 -7914 523 -7897
rect 755 -7914 772 -7897
rect 921 -7914 938 -7897
rect 423 -7914 440 -7897
rect 672 -8148 689 -8131
rect 506 -8148 523 -8131
rect 755 -8148 772 -8131
rect 921 -8148 938 -8131
rect 257 -8148 274 -8131
rect 672 -8382 689 -8365
rect 506 -8382 523 -8365
rect 755 -8382 772 -8365
rect 921 -8382 938 -8365
rect 257 -8382 274 -8365
rect 423 -8382 440 -8365
rect 174 -8616 191 -8599
rect 672 -8616 689 -8599
rect 755 -8616 772 -8599
rect 506 -8616 523 -8599
rect 921 -8616 938 -8599
rect 174 -8850 191 -8833
rect 672 -8850 689 -8833
rect 755 -8850 772 -8833
rect 506 -8850 523 -8833
rect 921 -8850 938 -8833
rect 423 -8850 440 -8833
rect 174 -9084 191 -9067
rect 672 -9084 689 -9067
rect 755 -9084 772 -9067
rect 506 -9084 523 -9067
rect 921 -9084 938 -9067
rect 257 -9084 274 -9067
rect 174 -9318 191 -9301
rect 672 -9318 689 -9301
rect 755 -9318 772 -9301
rect 506 -9318 523 -9301
rect 921 -9318 938 -9301
rect 257 -9318 274 -9301
rect 423 -9318 440 -9301
rect 672 -9552 689 -9535
rect 506 -9552 523 -9535
rect 755 -9552 772 -9535
rect 921 -9552 938 -9535
rect 8 -9552 25 -9535
rect 672 -9786 689 -9769
rect 506 -9786 523 -9769
rect 755 -9786 772 -9769
rect 921 -9786 938 -9769
rect 8 -9786 25 -9769
rect 423 -9786 440 -9769
rect 672 -10020 689 -10003
rect 506 -10020 523 -10003
rect 755 -10020 772 -10003
rect 921 -10020 938 -10003
rect 257 -10020 274 -10003
rect 8 -10020 25 -10003
rect 672 -10254 689 -10237
rect 506 -10254 523 -10237
rect 755 -10254 772 -10237
rect 921 -10254 938 -10237
rect 257 -10254 274 -10237
rect 8 -10254 25 -10237
rect 423 -10254 440 -10237
rect 174 -10488 191 -10471
rect 672 -10488 689 -10471
rect 755 -10488 772 -10471
rect 506 -10488 523 -10471
rect 921 -10488 938 -10471
rect 8 -10488 25 -10471
rect 174 -10722 191 -10705
rect 672 -10722 689 -10705
rect 755 -10722 772 -10705
rect 506 -10722 523 -10705
rect 921 -10722 938 -10705
rect 8 -10722 25 -10705
rect 423 -10722 440 -10705
rect 174 -10956 191 -10939
rect 672 -10956 689 -10939
rect 755 -10956 772 -10939
rect 506 -10956 523 -10939
rect 921 -10956 938 -10939
rect 257 -10956 274 -10939
rect 8 -10956 25 -10939
rect 174 -11190 191 -11173
rect 672 -11190 689 -11173
rect 755 -11190 772 -11173
rect 921 -11190 938 -11173
rect 257 -11190 274 -11173
rect 8 -11190 25 -11173
rect 423 -11190 440 -11173
rect 506 -11424 523 -11407
rect 755 -11424 772 -11407
rect 672 -11658 689 -11641
rect 921 -11658 938 -11641
rect 257 -11658 274 -11641
rect 423 -11658 440 -11641
rect 174 -11892 191 -11875
rect 672 -11892 689 -11875
rect 506 -11892 523 -11875
rect 755 -11892 772 -11875
rect 921 -11892 938 -11875
rect 257 -11892 274 -11875
rect 423 -11892 440 -11875
rect 174 -12126 191 -12109
rect 672 -12126 689 -12109
rect 755 -12126 772 -12109
rect 921 -12126 938 -12109
rect 257 -12126 274 -12109
rect 8 -12126 25 -12109
rect 506 -12360 523 -12343
rect 257 -12360 274 -12343
rect 8 -12360 25 -12343
rect 423 -12360 440 -12343
rect 174 -12594 191 -12577
rect 672 -12594 689 -12577
rect 755 -12594 772 -12577
rect 506 -12594 523 -12577
rect 8 -12594 25 -12577
rect 423 -12594 440 -12577
rect 174 -12828 191 -12811
rect 672 -12828 689 -12811
rect 506 -12828 523 -12811
rect 755 -12828 772 -12811
rect 921 -12828 938 -12811
rect 257 -12828 274 -12811
rect 8 -12828 25 -12811
rect 423 -12828 440 -12811
rect 174 -13062 191 -13045
rect 672 -13062 689 -13045
rect 506 -13062 523 -13045
rect 921 -13062 938 -13045
rect 755 -13062 772 -13045
rect 257 -13062 274 -13045
rect 8 -13062 25 -13045
rect 423 -13062 440 -13045
rect 174 -13296 191 -13279
rect 672 -13296 689 -13279
rect 506 -13296 523 -13279
rect 921 -13296 938 -13279
rect 257 -13296 274 -13279
rect 8 -13296 25 -13279
rect 423 -13296 440 -13279
rect 174 -13530 191 -13513
rect 506 -13530 523 -13513
rect 755 -13530 772 -13513
rect 257 -13530 274 -13513
rect 8 -13530 25 -13513
rect 423 -13530 440 -13513
rect 174 -13764 191 -13747
rect 672 -13764 689 -13747
rect 755 -13764 772 -13747
rect 257 -13764 274 -13747
rect 8 -13764 25 -13747
rect 423 -13764 440 -13747
rect 506 -13998 523 -13981
rect 8 -13998 25 -13981
rect 423 -13998 440 -13981
rect 174 -14232 191 -14215
rect 672 -14232 689 -14215
rect 755 -14232 772 -14215
rect 506 -14232 523 -14215
rect 921 -14232 938 -14215
rect 257 -14232 274 -14215
rect 672 -14466 689 -14449
rect 506 -14466 523 -14449
rect 921 -14466 938 -14449
rect 257 -14466 274 -14449
rect 423 -14466 440 -14449
rect 672 -14700 689 -14683
rect 506 -14700 523 -14683
rect 755 -14700 772 -14683
rect 921 -14700 938 -14683
rect 423 -14700 440 -14683
rect 755 -14934 772 -14917
<< poly >>
rect -51 -17 996 0
rect -51 -134 996 -117
rect -51 -251 996 -234
rect -51 -368 996 -351
rect -51 -485 996 -468
rect -51 -602 996 -585
rect -51 -719 996 -702
rect -51 -836 996 -819
rect -51 -953 996 -936
rect -51 -1070 996 -1053
rect -51 -1187 996 -1170
rect -51 -1304 996 -1287
rect -51 -1421 996 -1404
rect -51 -1538 996 -1521
rect -51 -1655 996 -1638
rect -51 -1772 996 -1755
rect -51 -1889 996 -1872
rect -51 -2006 996 -1989
rect -51 -2123 996 -2106
rect -51 -2240 996 -2223
rect -51 -2357 996 -2340
rect -51 -2474 996 -2457
rect -51 -2591 996 -2574
rect -51 -2708 996 -2691
rect -51 -2825 996 -2808
rect -51 -2942 996 -2925
rect -51 -3059 996 -3042
rect -51 -3176 996 -3159
rect -51 -3293 996 -3276
rect -51 -3410 996 -3393
rect -51 -3527 996 -3510
rect -51 -3644 996 -3627
rect -51 -3761 996 -3744
rect -51 -3878 996 -3861
rect -51 -3995 996 -3978
rect -51 -4112 996 -4095
rect -51 -4229 996 -4212
rect -51 -4346 996 -4329
rect -51 -4463 996 -4446
rect -51 -4580 996 -4563
rect -51 -4697 996 -4680
rect -51 -4814 996 -4797
rect -51 -4931 996 -4914
rect -51 -5048 996 -5031
rect -51 -5165 996 -5148
rect -51 -5282 996 -5265
rect -51 -5399 996 -5382
rect -51 -5516 996 -5499
rect -51 -5633 996 -5616
rect -51 -5750 996 -5733
rect -51 -5867 996 -5850
rect -51 -5984 996 -5967
rect -51 -6101 996 -6084
rect -51 -6218 996 -6201
rect -51 -6335 996 -6318
rect -51 -6452 996 -6435
rect -51 -6569 996 -6552
rect -51 -6686 996 -6669
rect -51 -6803 996 -6786
rect -51 -6920 996 -6903
rect -51 -7037 996 -7020
rect -51 -7154 996 -7137
rect -51 -7271 996 -7254
rect -51 -7388 996 -7371
rect -51 -7505 996 -7488
rect -51 -7622 996 -7605
rect -51 -7739 996 -7722
rect -51 -7856 996 -7839
rect -51 -7973 996 -7956
rect -51 -8090 996 -8073
rect -51 -8207 996 -8190
rect -51 -8324 996 -8307
rect -51 -8441 996 -8424
rect -51 -8558 996 -8541
rect -51 -8675 996 -8658
rect -51 -8792 996 -8775
rect -51 -8909 996 -8892
rect -51 -9026 996 -9009
rect -51 -9143 996 -9126
rect -51 -9260 996 -9243
rect -51 -9377 996 -9360
rect -51 -9494 996 -9477
rect -51 -9611 996 -9594
rect -51 -9728 996 -9711
rect -51 -9845 996 -9828
rect -51 -9962 996 -9945
rect -51 -10079 996 -10062
rect -51 -10196 996 -10179
rect -51 -10313 996 -10296
rect -51 -10430 996 -10413
rect -51 -10547 996 -10530
rect -51 -10664 996 -10647
rect -51 -10781 996 -10764
rect -51 -10898 996 -10881
rect -51 -11015 996 -10998
rect -51 -11132 996 -11115
rect -51 -11249 996 -11232
rect -51 -11366 996 -11349
rect -51 -11483 996 -11466
rect -51 -11600 996 -11583
rect -51 -11717 996 -11700
rect -51 -11834 996 -11817
rect -51 -11951 996 -11934
rect -51 -12068 996 -12051
rect -51 -12185 996 -12168
rect -51 -12302 996 -12285
rect -51 -12419 996 -12402
rect -51 -12536 996 -12519
rect -51 -12653 996 -12636
rect -51 -12770 996 -12753
rect -51 -12887 996 -12870
rect -51 -13004 996 -12987
rect -51 -13121 996 -13104
rect -51 -13238 996 -13221
rect -51 -13355 996 -13338
rect -51 -13472 996 -13455
rect -51 -13589 996 -13572
rect -51 -13706 996 -13689
rect -51 -13823 996 -13806
rect -51 -13940 996 -13923
rect -51 -14057 996 -14040
rect -51 -14174 996 -14157
rect -51 -14291 996 -14274
rect -51 -14408 996 -14391
rect -51 -14525 996 -14508
rect -51 -14642 996 -14625
rect -51 -14759 996 -14742
rect -51 -14876 996 -14859
rect -60 166 -27 199
rect -27 174 986 191
<< polycont >>
rect -52 174 -35 191
<< locali >>
rect 0 -14976 33 41
rect 83 -14976 116 41
rect 166 -14976 199 41
rect 249 -14976 282 41
rect 332 -14976 365 41
rect 415 -14976 448 41
rect 498 -14976 531 41
rect 581 -14976 614 41
rect 664 -14976 697 41
rect 747 -14976 780 41
rect 830 -14976 863 41
rect 913 -14976 946 41
rect 913 19 946 52
rect 913 138 946 171
rect 904 194 955 227
rect 904 227 955 244
rect 747 19 780 52
rect 747 138 780 171
rect 738 194 789 227
rect 738 227 789 244
rect 664 19 697 52
rect 664 138 697 171
rect 655 194 706 227
rect 655 227 706 244
rect 498 19 531 52
rect 498 138 531 171
rect 489 194 540 227
rect 489 227 540 244
rect 415 19 448 52
rect 415 138 448 171
rect 406 194 457 227
rect 406 227 457 244
rect 249 19 282 52
rect 249 138 282 171
rect 240 194 291 227
rect 240 227 291 244
rect 166 19 199 52
rect 166 138 199 171
rect 157 194 208 227
rect 157 227 208 244
rect 0 19 33 52
rect 0 138 33 171
rect -9 194 42 227
rect -9 227 42 244
rect -27 69 973 117
rect -60 69 -27 199
rect 830 41 863 69
rect 581 41 614 69
rect 332 41 365 69
rect 83 41 116 69
rect -25 244 971 292
<< viali >>
rect 921 27 938 44
rect 921 146 938 163
rect 755 27 772 44
rect 755 146 772 163
rect 672 27 689 44
rect 672 146 689 163
rect 506 27 523 44
rect 506 146 523 163
rect 423 27 440 44
rect 423 146 440 163
rect 257 27 274 44
rect 257 146 274 163
rect 174 27 191 44
rect 174 146 191 163
rect 8 27 25 44
rect 8 146 25 163
<< metal1 >>
rect 913 19 946 171
rect 747 19 780 171
rect 664 19 697 171
rect 498 19 531 171
rect 415 19 448 171
rect 249 19 282 171
rect 166 19 199 171
rect 0 19 33 171
<< end >>