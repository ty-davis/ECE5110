magic
tech sky130A
timestamp 1741801383
<< nwell >>
rect 11 197 314 488
<< nmos >>
rect 81 113 96 163
rect 135 113 150 163
rect 171 113 186 163
rect 224 113 239 163
<< pmos >>
rect 90 315 105 415
rect 126 315 141 415
rect 180 315 195 415
rect 216 315 231 415
<< ndiff >>
rect 45 155 81 163
rect 45 121 53 155
rect 70 121 81 155
rect 45 113 81 121
rect 96 155 135 163
rect 96 121 107 155
rect 124 121 135 155
rect 96 113 135 121
rect 150 113 171 163
rect 186 155 224 163
rect 186 121 196 155
rect 213 121 224 155
rect 186 113 224 121
rect 239 155 275 163
rect 239 121 250 155
rect 267 121 275 155
rect 239 113 275 121
<< pdiff >>
rect 54 407 90 415
rect 54 323 62 407
rect 79 323 90 407
rect 54 315 90 323
rect 105 315 126 415
rect 141 407 180 415
rect 141 323 152 407
rect 169 323 180 407
rect 141 315 180 323
rect 195 315 216 415
rect 231 407 267 415
rect 231 323 242 407
rect 259 323 267 407
rect 231 315 267 323
<< ndiffc >>
rect 53 121 70 155
rect 107 121 124 155
rect 196 121 213 155
rect 250 121 267 155
<< pdiffc >>
rect 62 323 79 407
rect 152 323 169 407
rect 242 323 259 407
<< psubdiff >>
rect 13 10 25 38
rect 300 10 312 38
<< nsubdiff >>
rect 29 442 41 470
rect 284 442 296 470
<< psubdiffcont >>
rect 25 10 300 38
<< nsubdiffcont >>
rect 41 442 284 470
<< poly >>
rect 90 415 105 428
rect 126 415 141 428
rect 180 415 195 428
rect 216 415 231 428
rect 90 298 105 315
rect 54 290 105 298
rect 54 273 62 290
rect 79 276 105 290
rect 79 273 87 276
rect 54 265 87 273
rect 72 194 87 265
rect 126 252 141 315
rect 180 252 195 315
rect 216 297 231 315
rect 216 289 282 297
rect 216 281 257 289
rect 108 244 141 252
rect 108 227 116 244
rect 133 227 141 244
rect 108 219 141 227
rect 162 244 195 252
rect 162 227 170 244
rect 187 227 195 244
rect 162 219 195 227
rect 126 195 141 219
rect 180 195 195 219
rect 72 179 96 194
rect 126 180 150 195
rect 81 163 96 179
rect 135 163 150 180
rect 171 180 195 195
rect 234 272 257 281
rect 274 272 282 289
rect 234 264 282 272
rect 234 186 249 264
rect 171 163 186 180
rect 224 171 249 186
rect 224 163 239 171
rect 81 100 96 113
rect 135 100 150 113
rect 171 100 186 113
rect 224 100 239 113
<< polycont >>
rect 62 273 79 290
rect 116 227 133 244
rect 170 227 187 244
rect 257 272 274 289
<< locali >>
rect 13 470 312 480
rect 13 442 41 470
rect 284 442 312 470
rect 13 432 312 442
rect 54 407 87 432
rect 54 323 62 407
rect 79 323 87 407
rect 54 315 87 323
rect 144 407 177 415
rect 144 323 152 407
rect 169 323 177 407
rect 54 290 87 298
rect 54 273 62 290
rect 79 273 87 290
rect 54 265 87 273
rect 144 288 177 323
rect 234 407 267 432
rect 234 323 242 407
rect 259 323 267 407
rect 234 315 267 323
rect 249 289 282 297
rect 144 271 231 288
rect 108 244 141 252
rect 108 227 116 244
rect 133 227 141 244
rect 108 219 141 227
rect 162 244 195 252
rect 162 227 170 244
rect 187 227 195 244
rect 162 219 195 227
rect 212 228 231 271
rect 249 272 257 289
rect 274 272 282 289
rect 249 264 282 272
rect 249 228 282 239
rect 212 206 282 228
rect 212 203 231 206
rect 45 180 169 200
rect 45 155 78 180
rect 45 121 53 155
rect 70 121 78 155
rect 45 113 78 121
rect 99 155 132 163
rect 99 121 107 155
rect 124 121 132 155
rect 99 48 132 121
rect 152 84 169 180
rect 202 186 231 203
rect 202 168 221 186
rect 188 155 221 168
rect 188 121 196 155
rect 213 121 221 155
rect 188 113 221 121
rect 242 155 275 163
rect 242 121 250 155
rect 267 121 275 155
rect 242 84 275 121
rect 152 67 275 84
rect 13 38 312 48
rect 13 10 25 38
rect 300 10 312 38
rect 13 0 312 10
<< labels >>
flabel pdiff 195 365 195 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 126 363 126 363 1 FreeSerif 8 0 0 0 S$
flabel pdiff 231 365 231 365 1 FreeSerif 8 0 0 0 S$
flabel pdiff 90 365 90 365 1 FreeSerif 8 0 0 0 S$
flabel locali 249 264 282 297 0 FreeSerif 80 0 0 0 B
port 14 nsew
flabel ndiff 135 137 135 137 1 FreeSerif 8 0 0 0 S$
flabel ndiff 171 137 171 137 1 FreeSerif 8 0 0 0 S$
flabel ndiff 96 135 96 135 1 FreeSerif 8 0 0 0 S$
flabel ndiff 239 138 239 138 1 FreeSerif 8 0 0 0 S$
flabel locali 162 219 195 252 0 FreeSerif 80 0 0 0 ~A
port 13 nsew
flabel locali 54 265 87 298 0 FreeSerif 80 0 0 0 A
port 11 nsew
flabel locali 108 219 141 252 0 FreeSerif 80 0 0 0 ~B
port 12 nsew
flabel locali 249 206 282 239 0 FreeSerif 80 0 0 0 Y
port 4 nsew
flabel locali 13 432 312 480 0 FreeSerif 80 0 0 0 VDD!
port 2 nsew
flabel locali 13 0 312 48 0 FreeSerif 80 0 0 0 GND!
port 3 nsew
<< end >>
